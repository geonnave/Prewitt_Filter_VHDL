library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.filter_masks.all;

package max_constants is
	constant	MMLength	:	integer	:=	25;
end;
