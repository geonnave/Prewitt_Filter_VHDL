library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.mem_size.all;
use work.matrix_types.all;

entity MemImgROM is
	port
	(
		addr_i	:	in	natural		range 0 to lin;
		addr_j	:	in	natural		range 0 to col;
		clk		:	in std_logic;
		q		:	out matrix_in
	);
end entity;


architecture rtl of MemImgROM is

	-- Build a 2-D array type for the RoM
	subtype pixel is std_logic_vector(7 downto 0);
	type memory_t is array(0 to lin, 0 to col) of pixel;
		
	function init_rom
		return memory_t is
		variable tmp : memory_t;
		begin
			tmp(0,0) := "00000000";
			tmp(41,0) := "00000000";
			tmp(0,1) := "00000000";
			tmp(41,1) := "00000000";
			tmp(0,2) := "00000000";
			tmp(41,2) := "00000000";
			tmp(0,3) := "00000000";
			tmp(41,3) := "00000000";
			tmp(0,4) := "00000000";
			tmp(41,4) := "00000000";
			tmp(0,5) := "00000000";
			tmp(41,5) := "00000000";
			tmp(0,6) := "00000000";
			tmp(41,6) := "00000000";
			tmp(0,7) := "00000000";
			tmp(41,7) := "00000000";
			tmp(0,8) := "00000000";
			tmp(41,8) := "00000000";
			tmp(0,9) := "00000000";
			tmp(41,9) := "00000000";
			tmp(0,10) := "00000000";
			tmp(41,10) := "00000000";
			tmp(0,11) := "00000000";
			tmp(41,11) := "00000000";
			tmp(0,12) := "00000000";
			tmp(41,12) := "00000000";
			tmp(0,13) := "00000000";
			tmp(41,13) := "00000000";
			tmp(0,14) := "00000000";
			tmp(41,14) := "00000000";
			tmp(0,15) := "00000000";
			tmp(41,15) := "00000000";
			tmp(0,16) := "00000000";
			tmp(41,16) := "00000000";
			tmp(0,17) := "00000000";
			tmp(41,17) := "00000000";
			tmp(0,18) := "00000000";
			tmp(41,18) := "00000000";
			tmp(0,19) := "00000000";
			tmp(41,19) := "00000000";
			tmp(0,20) := "00000000";
			tmp(41,20) := "00000000";
			tmp(0,21) := "00000000";
			tmp(41,21) := "00000000";
			tmp(0,22) := "00000000";
			tmp(41,22) := "00000000";
			tmp(0,23) := "00000000";
			tmp(41,23) := "00000000";
			tmp(0,24) := "00000000";
			tmp(41,24) := "00000000";
			tmp(0,25) := "00000000";
			tmp(41,25) := "00000000";
			tmp(0,26) := "00000000";
			tmp(41,26) := "00000000";
			tmp(0,27) := "00000000";
			tmp(41,27) := "00000000";
			tmp(0,28) := "00000000";
			tmp(41,28) := "00000000";
			tmp(0,29) := "00000000";
			tmp(41,29) := "00000000";
			tmp(0,30) := "00000000";
			tmp(41,30) := "00000000";
			tmp(0,31) := "00000000";
			tmp(41,31) := "00000000";
			tmp(0,32) := "00000000";
			tmp(41,32) := "00000000";
			tmp(0,33) := "00000000";
			tmp(41,33) := "00000000";
			tmp(0,34) := "00000000";
			tmp(41,34) := "00000000";
			tmp(0,35) := "00000000";
			tmp(41,35) := "00000000";
			tmp(0,36) := "00000000";
			tmp(41,36) := "00000000";
			tmp(0,37) := "00000000";
			tmp(41,37) := "00000000";
			tmp(0,38) := "00000000";
			tmp(41,38) := "00000000";
			tmp(0,39) := "00000000";
			tmp(41,39) := "00000000";
			tmp(0,40) := "00000000";
			tmp(41,40) := "00000000";
			tmp(0,41) := "00000000";
			tmp(41,41) := "00000000";
			tmp(0,0) := "00000000";
			tmp(0,41) := "00000000";
			tmp(1,0) := "00000000";
			tmp(1,41) := "00000000";
			tmp(2,0) := "00000000";
			tmp(2,41) := "00000000";
			tmp(3,0) := "00000000";
			tmp(3,41) := "00000000";
			tmp(4,0) := "00000000";
			tmp(4,41) := "00000000";
			tmp(5,0) := "00000000";
			tmp(5,41) := "00000000";
			tmp(6,0) := "00000000";
			tmp(6,41) := "00000000";
			tmp(7,0) := "00000000";
			tmp(7,41) := "00000000";
			tmp(8,0) := "00000000";
			tmp(8,41) := "00000000";
			tmp(9,0) := "00000000";
			tmp(9,41) := "00000000";
			tmp(10,0) := "00000000";
			tmp(10,41) := "00000000";
			tmp(11,0) := "00000000";
			tmp(11,41) := "00000000";
			tmp(12,0) := "00000000";
			tmp(12,41) := "00000000";
			tmp(13,0) := "00000000";
			tmp(13,41) := "00000000";
			tmp(14,0) := "00000000";
			tmp(14,41) := "00000000";
			tmp(15,0) := "00000000";
			tmp(15,41) := "00000000";
			tmp(16,0) := "00000000";
			tmp(16,41) := "00000000";
			tmp(17,0) := "00000000";
			tmp(17,41) := "00000000";
			tmp(18,0) := "00000000";
			tmp(18,41) := "00000000";
			tmp(19,0) := "00000000";
			tmp(19,41) := "00000000";
			tmp(20,0) := "00000000";
			tmp(20,41) := "00000000";
			tmp(21,0) := "00000000";
			tmp(21,41) := "00000000";
			tmp(22,0) := "00000000";
			tmp(22,41) := "00000000";
			tmp(23,0) := "00000000";
			tmp(23,41) := "00000000";
			tmp(24,0) := "00000000";
			tmp(24,41) := "00000000";
			tmp(25,0) := "00000000";
			tmp(25,41) := "00000000";
			tmp(26,0) := "00000000";
			tmp(26,41) := "00000000";
			tmp(27,0) := "00000000";
			tmp(27,41) := "00000000";
			tmp(28,0) := "00000000";
			tmp(28,41) := "00000000";
			tmp(29,0) := "00000000";
			tmp(29,41) := "00000000";
			tmp(30,0) := "00000000";
			tmp(30,41) := "00000000";
			tmp(31,0) := "00000000";
			tmp(31,41) := "00000000";
			tmp(32,0) := "00000000";
			tmp(32,41) := "00000000";
			tmp(33,0) := "00000000";
			tmp(33,41) := "00000000";
			tmp(34,0) := "00000000";
			tmp(34,41) := "00000000";
			tmp(35,0) := "00000000";
			tmp(35,41) := "00000000";
			tmp(36,0) := "00000000";
			tmp(36,41) := "00000000";
			tmp(37,0) := "00000000";
			tmp(37,41) := "00000000";
			tmp(38,0) := "00000000";
			tmp(38,41) := "00000000";
			tmp(39,0) := "00000000";
			tmp(39,41) := "00000000";
			tmp(40,0) := "00000000";
			tmp(40,41) := "00000000";
			tmp(41,0) := "00000000";
			tmp(41,41) := "00000000";
			tmp(1,1) := "10100001";
			tmp(1,2) := "00100001";
			tmp(1,3) := "00000000";
			tmp(1,4) := "00000000";
			tmp(1,5) := "00011000";
			tmp(1,6) := "11001101";
			tmp(1,7) := "11111110";
			tmp(1,8) := "11111111";
			tmp(1,9) := "11111100";
			tmp(1,10) := "11011000";
			tmp(1,11) := "01000001";
			tmp(1,12) := "00000000";
			tmp(1,13) := "00000010";
			tmp(1,14) := "00001101";
			tmp(1,15) := "00000000";
			tmp(1,16) := "00100010";
			tmp(1,17) := "01101010";
			tmp(1,18) := "10001010";
			tmp(1,19) := "01001001";
			tmp(1,20) := "00101100";
			tmp(1,21) := "00010100";
			tmp(1,22) := "00000010";
			tmp(1,23) := "00000001";
			tmp(1,24) := "00100101";
			tmp(1,25) := "10110101";
			tmp(1,26) := "11111000";
			tmp(1,27) := "11110101";
			tmp(1,28) := "11110110";
			tmp(1,29) := "11111000";
			tmp(1,30) := "11110111";
			tmp(1,31) := "11110011";
			tmp(1,32) := "11100011";
			tmp(1,33) := "10110011";
			tmp(1,34) := "01111101";
			tmp(1,35) := "01100000";
			tmp(1,36) := "01011101";
			tmp(1,37) := "01011000";
			tmp(1,38) := "01010101";
			tmp(1,39) := "01010100";
			tmp(1,40) := "01010010";
			tmp(2,1) := "10110001";
			tmp(2,2) := "00011000";
			tmp(2,3) := "00000000";
			tmp(2,4) := "00000000";
			tmp(2,5) := "00100010";
			tmp(2,6) := "11001001";
			tmp(2,7) := "11111101";
			tmp(2,8) := "11111111";
			tmp(2,9) := "11111010";
			tmp(2,10) := "11010101";
			tmp(2,11) := "01001101";
			tmp(2,12) := "00010010";
			tmp(2,13) := "00011100";
			tmp(2,14) := "01011010";
			tmp(2,15) := "10010101";
			tmp(2,16) := "10110011";
			tmp(2,17) := "01110110";
			tmp(2,18) := "00001010";
			tmp(2,19) := "00001100";
			tmp(2,20) := "00000000";
			tmp(2,21) := "00000000";
			tmp(2,22) := "00000000";
			tmp(2,23) := "00000000";
			tmp(2,24) := "00100001";
			tmp(2,25) := "10110000";
			tmp(2,26) := "11110101";
			tmp(2,27) := "11110110";
			tmp(2,28) := "11111010";
			tmp(2,29) := "11111001";
			tmp(2,30) := "11100110";
			tmp(2,31) := "11000101";
			tmp(2,32) := "10101001";
			tmp(2,33) := "10001001";
			tmp(2,34) := "01101100";
			tmp(2,35) := "01100011";
			tmp(2,36) := "01011110";
			tmp(2,37) := "01011100";
			tmp(2,38) := "01011000";
			tmp(2,39) := "01010111";
			tmp(2,40) := "01010110";
			tmp(3,1) := "10101100";
			tmp(3,2) := "00100010";
			tmp(3,3) := "00000111";
			tmp(3,4) := "00000000";
			tmp(3,5) := "00011111";
			tmp(3,6) := "10111100";
			tmp(3,7) := "11111100";
			tmp(3,8) := "11111101";
			tmp(3,9) := "11110000";
			tmp(3,10) := "11011001";
			tmp(3,11) := "01111001";
			tmp(3,12) := "10011011";
			tmp(3,13) := "11001000";
			tmp(3,14) := "11100101";
			tmp(3,15) := "11110111";
			tmp(3,16) := "11101111";
			tmp(3,17) := "10001110";
			tmp(3,18) := "00001101";
			tmp(3,19) := "00000000";
			tmp(3,20) := "00000000";
			tmp(3,21) := "00000000";
			tmp(3,22) := "00000110";
			tmp(3,23) := "00000111";
			tmp(3,24) := "00100000";
			tmp(3,25) := "10101101";
			tmp(3,26) := "11110110";
			tmp(3,27) := "11111010";
			tmp(3,28) := "11110000";
			tmp(3,29) := "11011111";
			tmp(3,30) := "10111111";
			tmp(3,31) := "10010100";
			tmp(3,32) := "01110111";
			tmp(3,33) := "01101011";
			tmp(3,34) := "01100110";
			tmp(3,35) := "01100101";
			tmp(3,36) := "01100001";
			tmp(3,37) := "01011110";
			tmp(3,38) := "01011100";
			tmp(3,39) := "01011011";
			tmp(3,40) := "01011011";
			tmp(4,1) := "10101100";
			tmp(4,2) := "00100110";
			tmp(4,3) := "00000000";
			tmp(4,4) := "00000001";
			tmp(4,5) := "00101110";
			tmp(4,6) := "10111001";
			tmp(4,7) := "11101100";
			tmp(4,8) := "10111100";
			tmp(4,9) := "01111000";
			tmp(4,10) := "01010010";
			tmp(4,11) := "11000001";
			tmp(4,12) := "11110011";
			tmp(4,13) := "11111111";
			tmp(4,14) := "11111011";
			tmp(4,15) := "11111111";
			tmp(4,16) := "11111101";
			tmp(4,17) := "10010111";
			tmp(4,18) := "00001110";
			tmp(4,19) := "00000110";
			tmp(4,20) := "00000000";
			tmp(4,21) := "00000000";
			tmp(4,22) := "00000010";
			tmp(4,23) := "00000000";
			tmp(4,24) := "00010100";
			tmp(4,25) := "10100100";
			tmp(4,26) := "11110010";
			tmp(4,27) := "11110101";
			tmp(4,28) := "11010001";
			tmp(4,29) := "10101100";
			tmp(4,30) := "10010010";
			tmp(4,31) := "01111100";
			tmp(4,32) := "01110001";
			tmp(4,33) := "01110000";
			tmp(4,34) := "01110001";
			tmp(4,35) := "01100111";
			tmp(4,36) := "01100100";
			tmp(4,37) := "01100001";
			tmp(4,38) := "01011111";
			tmp(4,39) := "01011111";
			tmp(4,40) := "01011110";
			tmp(5,1) := "10101011";
			tmp(5,2) := "00100000";
			tmp(5,3) := "00001101";
			tmp(5,4) := "00101011";
			tmp(5,5) := "01100001";
			tmp(5,6) := "01100011";
			tmp(5,7) := "00111010";
			tmp(5,8) := "00001010";
			tmp(5,9) := "00001100";
			tmp(5,10) := "00110000";
			tmp(5,11) := "10101101";
			tmp(5,12) := "11110100";
			tmp(5,13) := "11111111";
			tmp(5,14) := "11110101";
			tmp(5,15) := "11111101";
			tmp(5,16) := "11101010";
			tmp(5,17) := "10010000";
			tmp(5,18) := "00010100";
			tmp(5,19) := "00000010";
			tmp(5,20) := "00000000";
			tmp(5,21) := "00000000";
			tmp(5,22) := "00000001";
			tmp(5,23) := "00000000";
			tmp(5,24) := "00011001";
			tmp(5,25) := "10101001";
			tmp(5,26) := "11110011";
			tmp(5,27) := "11011000";
			tmp(5,28) := "10101110";
			tmp(5,29) := "10001010";
			tmp(5,30) := "01111111";
			tmp(5,31) := "01111100";
			tmp(5,32) := "01111011";
			tmp(5,33) := "01111001";
			tmp(5,34) := "01110110";
			tmp(5,35) := "01101001";
			tmp(5,36) := "01100110";
			tmp(5,37) := "01100011";
			tmp(5,38) := "01100001";
			tmp(5,39) := "01100000";
			tmp(5,40) := "01100000";
			tmp(6,1) := "10101001";
			tmp(6,2) := "10000110";
			tmp(6,3) := "10111010";
			tmp(6,4) := "11010001";
			tmp(6,5) := "11001100";
			tmp(6,6) := "01001100";
			tmp(6,7) := "00000111";
			tmp(6,8) := "00000000";
			tmp(6,9) := "00000100";
			tmp(6,10) := "00010101";
			tmp(6,11) := "10101011";
			tmp(6,12) := "11110101";
			tmp(6,13) := "11111110";
			tmp(6,14) := "11111111";
			tmp(6,15) := "11111111";
			tmp(6,16) := "11110100";
			tmp(6,17) := "10011001";
			tmp(6,18) := "00010001";
			tmp(6,19) := "00000011";
			tmp(6,20) := "00000001";
			tmp(6,21) := "00000101";
			tmp(6,22) := "00000100";
			tmp(6,23) := "00000101";
			tmp(6,24) := "00011111";
			tmp(6,25) := "10011110";
			tmp(6,26) := "11010100";
			tmp(6,27) := "10110000";
			tmp(6,28) := "10011000";
			tmp(6,29) := "10001000";
			tmp(6,30) := "10000100";
			tmp(6,31) := "01111111";
			tmp(6,32) := "01111001";
			tmp(6,33) := "01110100";
			tmp(6,34) := "01101110";
			tmp(6,35) := "01101011";
			tmp(6,36) := "01101001";
			tmp(6,37) := "01100101";
			tmp(6,38) := "01100011";
			tmp(6,39) := "01100010";
			tmp(6,40) := "01100001";
			tmp(7,1) := "01101001";
			tmp(7,2) := "11010100";
			tmp(7,3) := "11110010";
			tmp(7,4) := "11111111";
			tmp(7,5) := "11110111";
			tmp(7,6) := "01001011";
			tmp(7,7) := "00001000";
			tmp(7,8) := "00000110";
			tmp(7,9) := "00001000";
			tmp(7,10) := "00010011";
			tmp(7,11) := "10101110";
			tmp(7,12) := "11111100";
			tmp(7,13) := "11111111";
			tmp(7,14) := "11111101";
			tmp(7,15) := "11111111";
			tmp(7,16) := "11110000";
			tmp(7,17) := "10100000";
			tmp(7,18) := "00001101";
			tmp(7,19) := "00000000";
			tmp(7,20) := "00000000";
			tmp(7,21) := "00000001";
			tmp(7,22) := "00000000";
			tmp(7,23) := "00000000";
			tmp(7,24) := "00011000";
			tmp(7,25) := "10000100";
			tmp(7,26) := "10100001";
			tmp(7,27) := "10011001";
			tmp(7,28) := "10010000";
			tmp(7,29) := "10001011";
			tmp(7,30) := "10000110";
			tmp(7,31) := "01111100";
			tmp(7,32) := "01110110";
			tmp(7,33) := "01110011";
			tmp(7,34) := "01101100";
			tmp(7,35) := "01110000";
			tmp(7,36) := "01101101";
			tmp(7,37) := "01101001";
			tmp(7,38) := "01100110";
			tmp(7,39) := "01100110";
			tmp(7,40) := "01100011";
			tmp(8,1) := "01000111";
			tmp(8,2) := "11011001";
			tmp(8,3) := "11111111";
			tmp(8,4) := "11111111";
			tmp(8,5) := "11110011";
			tmp(8,6) := "01000111";
			tmp(8,7) := "00001000";
			tmp(8,8) := "00000000";
			tmp(8,9) := "00000000";
			tmp(8,10) := "00100000";
			tmp(8,11) := "10100011";
			tmp(8,12) := "11110110";
			tmp(8,13) := "11111101";
			tmp(8,14) := "11110110";
			tmp(8,15) := "11111011";
			tmp(8,16) := "11110100";
			tmp(8,17) := "10101110";
			tmp(8,18) := "00010010";
			tmp(8,19) := "00000000";
			tmp(8,20) := "00000001";
			tmp(8,21) := "00000100";
			tmp(8,22) := "00000000";
			tmp(8,23) := "00001001";
			tmp(8,24) := "00101001";
			tmp(8,25) := "10010000";
			tmp(8,26) := "10100011";
			tmp(8,27) := "10010111";
			tmp(8,28) := "10001110";
			tmp(8,29) := "10000110";
			tmp(8,30) := "01111110";
			tmp(8,31) := "01111001";
			tmp(8,32) := "01111100";
			tmp(8,33) := "01111011";
			tmp(8,34) := "01110011";
			tmp(8,35) := "01110011";
			tmp(8,36) := "01110000";
			tmp(8,37) := "01101011";
			tmp(8,38) := "01101000";
			tmp(8,39) := "01100111";
			tmp(8,40) := "01100101";
			tmp(9,1) := "00111101";
			tmp(9,2) := "11010001";
			tmp(9,3) := "11111100";
			tmp(9,4) := "11111111";
			tmp(9,5) := "11101100";
			tmp(9,6) := "01011011";
			tmp(9,7) := "00000000";
			tmp(9,8) := "00000101";
			tmp(9,9) := "00000010";
			tmp(9,10) := "00010110";
			tmp(9,11) := "10011101";
			tmp(9,12) := "11110111";
			tmp(9,13) := "11111111";
			tmp(9,14) := "11111100";
			tmp(9,15) := "11111101";
			tmp(9,16) := "11110110";
			tmp(9,17) := "10110001";
			tmp(9,18) := "00010010";
			tmp(9,19) := "00000101";
			tmp(9,20) := "00000001";
			tmp(9,21) := "00001001";
			tmp(9,22) := "00000000";
			tmp(9,23) := "00011101";
			tmp(9,24) := "01111010";
			tmp(9,25) := "10010111";
			tmp(9,26) := "10011100";
			tmp(9,27) := "10010011";
			tmp(9,28) := "10001101";
			tmp(9,29) := "10000101";
			tmp(9,30) := "10000001";
			tmp(9,31) := "01111110";
			tmp(9,32) := "01111100";
			tmp(9,33) := "01111010";
			tmp(9,34) := "01110110";
			tmp(9,35) := "01110001";
			tmp(9,36) := "01101111";
			tmp(9,37) := "01101101";
			tmp(9,38) := "01101000";
			tmp(9,39) := "01100111";
			tmp(9,40) := "01100101";
			tmp(10,1) := "00111101";
			tmp(10,2) := "11010001";
			tmp(10,3) := "11111100";
			tmp(10,4) := "11111111";
			tmp(10,5) := "11101101";
			tmp(10,6) := "01011110";
			tmp(10,7) := "00000000";
			tmp(10,8) := "00000101";
			tmp(10,9) := "00000010";
			tmp(10,10) := "00010110";
			tmp(10,11) := "10011011";
			tmp(10,12) := "11110110";
			tmp(10,13) := "11111111";
			tmp(10,14) := "11111011";
			tmp(10,15) := "11111110";
			tmp(10,16) := "11110111";
			tmp(10,17) := "10110010";
			tmp(10,18) := "00010011";
			tmp(10,19) := "00000000";
			tmp(10,20) := "00000001";
			tmp(10,21) := "00000000";
			tmp(10,22) := "00001000";
			tmp(10,23) := "01000111";
			tmp(10,24) := "10001100";
			tmp(10,25) := "10011100";
			tmp(10,26) := "10100010";
			tmp(10,27) := "10010010";
			tmp(10,28) := "10001101";
			tmp(10,29) := "10000101";
			tmp(10,30) := "10000001";
			tmp(10,31) := "01111111";
			tmp(10,32) := "01111110";
			tmp(10,33) := "01111010";
			tmp(10,34) := "01110111";
			tmp(10,35) := "01110010";
			tmp(10,36) := "01110000";
			tmp(10,37) := "01101101";
			tmp(10,38) := "01101010";
			tmp(10,39) := "01100111";
			tmp(10,40) := "01100101";
			tmp(11,1) := "00111101";
			tmp(11,2) := "11010001";
			tmp(11,3) := "11111100";
			tmp(11,4) := "11111111";
			tmp(11,5) := "11101111";
			tmp(11,6) := "01100010";
			tmp(11,7) := "00000000";
			tmp(11,8) := "00000100";
			tmp(11,9) := "00000001";
			tmp(11,10) := "00010100";
			tmp(11,11) := "10011000";
			tmp(11,12) := "11110101";
			tmp(11,13) := "11111111";
			tmp(11,14) := "11111011";
			tmp(11,15) := "11111110";
			tmp(11,16) := "11111001";
			tmp(11,17) := "10110101";
			tmp(11,18) := "00010110";
			tmp(11,19) := "00000000";
			tmp(11,20) := "00000011";
			tmp(11,21) := "00000000";
			tmp(11,22) := "00101110";
			tmp(11,23) := "01111100";
			tmp(11,24) := "10011011";
			tmp(11,25) := "10011110";
			tmp(11,26) := "10100001";
			tmp(11,27) := "10010010";
			tmp(11,28) := "10001100";
			tmp(11,29) := "10000101";
			tmp(11,30) := "10000001";
			tmp(11,31) := "10000000";
			tmp(11,32) := "01111110";
			tmp(11,33) := "01111010";
			tmp(11,34) := "01110111";
			tmp(11,35) := "01110100";
			tmp(11,36) := "01110010";
			tmp(11,37) := "01101111";
			tmp(11,38) := "01101011";
			tmp(11,39) := "01101001";
			tmp(11,40) := "01100110";
			tmp(12,1) := "00111000";
			tmp(12,2) := "11001110";
			tmp(12,3) := "11111110";
			tmp(12,4) := "11111111";
			tmp(12,5) := "11110010";
			tmp(12,6) := "01101000";
			tmp(12,7) := "00000000";
			tmp(12,8) := "00000011";
			tmp(12,9) := "00000001";
			tmp(12,10) := "00010010";
			tmp(12,11) := "10010100";
			tmp(12,12) := "11110100";
			tmp(12,13) := "11111111";
			tmp(12,14) := "11111011";
			tmp(12,15) := "11111110";
			tmp(12,16) := "11111011";
			tmp(12,17) := "10111010";
			tmp(12,18) := "00011001";
			tmp(12,19) := "00000010";
			tmp(12,20) := "00000100";
			tmp(12,21) := "00001010";
			tmp(12,22) := "01011100";
			tmp(12,23) := "10011010";
			tmp(12,24) := "10011010";
			tmp(12,25) := "10100010";
			tmp(12,26) := "10011000";
			tmp(12,27) := "10010000";
			tmp(12,28) := "10001011";
			tmp(12,29) := "10000101";
			tmp(12,30) := "10000010";
			tmp(12,31) := "10000001";
			tmp(12,32) := "01111111";
			tmp(12,33) := "01111011";
			tmp(12,34) := "01111000";
			tmp(12,35) := "01110110";
			tmp(12,36) := "01110100";
			tmp(12,37) := "01110000";
			tmp(12,38) := "01101101";
			tmp(12,39) := "01101010";
			tmp(12,40) := "01100111";
			tmp(13,1) := "00110100";
			tmp(13,2) := "11001001";
			tmp(13,3) := "11111101";
			tmp(13,4) := "11111111";
			tmp(13,5) := "11110101";
			tmp(13,6) := "01101110";
			tmp(13,7) := "00000001";
			tmp(13,8) := "00000011";
			tmp(13,9) := "00000001";
			tmp(13,10) := "00001111";
			tmp(13,11) := "10010000";
			tmp(13,12) := "11110001";
			tmp(13,13) := "11111111";
			tmp(13,14) := "11111010";
			tmp(13,15) := "11111110";
			tmp(13,16) := "11111101";
			tmp(13,17) := "10111100";
			tmp(13,18) := "00011101";
			tmp(13,19) := "00000100";
			tmp(13,20) := "00000001";
			tmp(13,21) := "00100110";
			tmp(13,22) := "10000010";
			tmp(13,23) := "10011100";
			tmp(13,24) := "10010100";
			tmp(13,25) := "10101000";
			tmp(13,26) := "10010001";
			tmp(13,27) := "10001111";
			tmp(13,28) := "10001011";
			tmp(13,29) := "10000110";
			tmp(13,30) := "10000011";
			tmp(13,31) := "10000010";
			tmp(13,32) := "10000000";
			tmp(13,33) := "01111101";
			tmp(13,34) := "01111001";
			tmp(13,35) := "01110111";
			tmp(13,36) := "01110110";
			tmp(13,37) := "01110010";
			tmp(13,38) := "01101110";
			tmp(13,39) := "01101010";
			tmp(13,40) := "01101000";
			tmp(14,1) := "00110000";
			tmp(14,2) := "11000110";
			tmp(14,3) := "11111110";
			tmp(14,4) := "11111101";
			tmp(14,5) := "11111000";
			tmp(14,6) := "01110100";
			tmp(14,7) := "00000011";
			tmp(14,8) := "00000010";
			tmp(14,9) := "00000000";
			tmp(14,10) := "00001101";
			tmp(14,11) := "10001011";
			tmp(14,12) := "11110001";
			tmp(14,13) := "11111111";
			tmp(14,14) := "11111010";
			tmp(14,15) := "11111110";
			tmp(14,16) := "11111111";
			tmp(14,17) := "11000000";
			tmp(14,18) := "00100001";
			tmp(14,19) := "00000000";
			tmp(14,20) := "00000101";
			tmp(14,21) := "01001010";
			tmp(14,22) := "10010110";
			tmp(14,23) := "10010100";
			tmp(14,24) := "10010100";
			tmp(14,25) := "10101011";
			tmp(14,26) := "10010011";
			tmp(14,27) := "10001110";
			tmp(14,28) := "10001010";
			tmp(14,29) := "10000101";
			tmp(14,30) := "10000011";
			tmp(14,31) := "10000011";
			tmp(14,32) := "10000010";
			tmp(14,33) := "01111110";
			tmp(14,34) := "01111010";
			tmp(14,35) := "01111000";
			tmp(14,36) := "01110110";
			tmp(14,37) := "01110010";
			tmp(14,38) := "01101110";
			tmp(14,39) := "01101011";
			tmp(14,40) := "01100111";
			tmp(15,1) := "00101111";
			tmp(15,2) := "11000110";
			tmp(15,3) := "11111110";
			tmp(15,4) := "11111011";
			tmp(15,5) := "11111010";
			tmp(15,6) := "01111000";
			tmp(15,7) := "00000101";
			tmp(15,8) := "00000001";
			tmp(15,9) := "00000000";
			tmp(15,10) := "00001100";
			tmp(15,11) := "10001000";
			tmp(15,12) := "11110000";
			tmp(15,13) := "11111111";
			tmp(15,14) := "11111001";
			tmp(15,15) := "11111110";
			tmp(15,16) := "11111111";
			tmp(15,17) := "11000010";
			tmp(15,18) := "00100011";
			tmp(15,19) := "00000000";
			tmp(15,20) := "00010100";
			tmp(15,21) := "01101100";
			tmp(15,22) := "10011010";
			tmp(15,23) := "10001111";
			tmp(15,24) := "10011100";
			tmp(15,25) := "10100100";
			tmp(15,26) := "10010110";
			tmp(15,27) := "10001101";
			tmp(15,28) := "10001001";
			tmp(15,29) := "10000101";
			tmp(15,30) := "10000100";
			tmp(15,31) := "10000100";
			tmp(15,32) := "10000010";
			tmp(15,33) := "01111110";
			tmp(15,34) := "01111011";
			tmp(15,35) := "01111000";
			tmp(15,36) := "01110110";
			tmp(15,37) := "01110010";
			tmp(15,38) := "01101110";
			tmp(15,39) := "01101010";
			tmp(15,40) := "01101000";
			tmp(16,1) := "00101111";
			tmp(16,2) := "11000110";
			tmp(16,3) := "11111101";
			tmp(16,4) := "11111100";
			tmp(16,5) := "11111011";
			tmp(16,6) := "01111011";
			tmp(16,7) := "00000101";
			tmp(16,8) := "00000001";
			tmp(16,9) := "00000000";
			tmp(16,10) := "00001011";
			tmp(16,11) := "10000110";
			tmp(16,12) := "11101111";
			tmp(16,13) := "11111111";
			tmp(16,14) := "11111001";
			tmp(16,15) := "11111110";
			tmp(16,16) := "11111111";
			tmp(16,17) := "11000100";
			tmp(16,18) := "00100101";
			tmp(16,19) := "00000000";
			tmp(16,20) := "00100110";
			tmp(16,21) := "10000011";
			tmp(16,22) := "10011001";
			tmp(16,23) := "10010010";
			tmp(16,24) := "10100100";
			tmp(16,25) := "10011010";
			tmp(16,26) := "10010110";
			tmp(16,27) := "10001100";
			tmp(16,28) := "10001001";
			tmp(16,29) := "10000101";
			tmp(16,30) := "10000100";
			tmp(16,31) := "10000101";
			tmp(16,32) := "10000011";
			tmp(16,33) := "01111111";
			tmp(16,34) := "01111011";
			tmp(16,35) := "01111000";
			tmp(16,36) := "01110101";
			tmp(16,37) := "01110010";
			tmp(16,38) := "01101110";
			tmp(16,39) := "01101010";
			tmp(16,40) := "01100110";
			tmp(17,1) := "00100001";
			tmp(17,2) := "11000101";
			tmp(17,3) := "11111111";
			tmp(17,4) := "11111111";
			tmp(17,5) := "11110001";
			tmp(17,6) := "10001010";
			tmp(17,7) := "00000000";
			tmp(17,8) := "00000110";
			tmp(17,9) := "00000000";
			tmp(17,10) := "00001011";
			tmp(17,11) := "10001000";
			tmp(17,12) := "11101010";
			tmp(17,13) := "11111111";
			tmp(17,14) := "11110111";
			tmp(17,15) := "11110101";
			tmp(17,16) := "11111111";
			tmp(17,17) := "11000100";
			tmp(17,18) := "00101010";
			tmp(17,19) := "00000000";
			tmp(17,20) := "00101011";
			tmp(17,21) := "10000101";
			tmp(17,22) := "10011101";
			tmp(17,23) := "10010000";
			tmp(17,24) := "10011111";
			tmp(17,25) := "10011010";
			tmp(17,26) := "10011000";
			tmp(17,27) := "10001011";
			tmp(17,28) := "10001000";
			tmp(17,29) := "10000101";
			tmp(17,30) := "10000100";
			tmp(17,31) := "10000010";
			tmp(17,32) := "01111111";
			tmp(17,33) := "01111100";
			tmp(17,34) := "01111010";
			tmp(17,35) := "01111001";
			tmp(17,36) := "01110110";
			tmp(17,37) := "01110010";
			tmp(17,38) := "01101111";
			tmp(17,39) := "01101101";
			tmp(17,40) := "01101010";
			tmp(18,1) := "00100010";
			tmp(18,2) := "10111000";
			tmp(18,3) := "11110000";
			tmp(18,4) := "11111110";
			tmp(18,5) := "11110001";
			tmp(18,6) := "10000111";
			tmp(18,7) := "00000001";
			tmp(18,8) := "00001101";
			tmp(18,9) := "00000010";
			tmp(18,10) := "00010001";
			tmp(18,11) := "01111100";
			tmp(18,12) := "11101110";
			tmp(18,13) := "11111110";
			tmp(18,14) := "11111110";
			tmp(18,15) := "11111111";
			tmp(18,16) := "11111111";
			tmp(18,17) := "11001101";
			tmp(18,18) := "00100011";
			tmp(18,19) := "00010000";
			tmp(18,20) := "01000100";
			tmp(18,21) := "10010110";
			tmp(18,22) := "10100000";
			tmp(18,23) := "10010011";
			tmp(18,24) := "10100011";
			tmp(18,25) := "10011010";
			tmp(18,26) := "10001100";
			tmp(18,27) := "10001011";
			tmp(18,28) := "10001000";
			tmp(18,29) := "10000101";
			tmp(18,30) := "10000011";
			tmp(18,31) := "10000010";
			tmp(18,32) := "10000001";
			tmp(18,33) := "01111100";
			tmp(18,34) := "01111010";
			tmp(18,35) := "01111000";
			tmp(18,36) := "01110101";
			tmp(18,37) := "01110010";
			tmp(18,38) := "01101111";
			tmp(18,39) := "01101101";
			tmp(18,40) := "01101010";
			tmp(19,1) := "00101111";
			tmp(19,2) := "10111101";
			tmp(19,3) := "11111001";
			tmp(19,4) := "11111111";
			tmp(19,5) := "11111010";
			tmp(19,6) := "10001010";
			tmp(19,7) := "00000000";
			tmp(19,8) := "00000000";
			tmp(19,9) := "00000000";
			tmp(19,10) := "00000111";
			tmp(19,11) := "01111001";
			tmp(19,12) := "11111100";
			tmp(19,13) := "11111000";
			tmp(19,14) := "11111111";
			tmp(19,15) := "11111111";
			tmp(19,16) := "11111010";
			tmp(19,17) := "11011101";
			tmp(19,18) := "00101010";
			tmp(19,19) := "00000000";
			tmp(19,20) := "01000001";
			tmp(19,21) := "10010010";
			tmp(19,22) := "10011001";
			tmp(19,23) := "10001101";
			tmp(19,24) := "10100000";
			tmp(19,25) := "10011101";
			tmp(19,26) := "10001111";
			tmp(19,27) := "10001011";
			tmp(19,28) := "10001000";
			tmp(19,29) := "10000101";
			tmp(19,30) := "10000011";
			tmp(19,31) := "10000010";
			tmp(19,32) := "10000000";
			tmp(19,33) := "01111101";
			tmp(19,34) := "01111010";
			tmp(19,35) := "01111000";
			tmp(19,36) := "01110101";
			tmp(19,37) := "01110001";
			tmp(19,38) := "01101110";
			tmp(19,39) := "01101100";
			tmp(19,40) := "01101001";
			tmp(20,1) := "00111100";
			tmp(20,2) := "10110010";
			tmp(20,3) := "11110101";
			tmp(20,4) := "11110010";
			tmp(20,5) := "11101000";
			tmp(20,6) := "10001110";
			tmp(20,7) := "00011110";
			tmp(20,8) := "00001010";
			tmp(20,9) := "00001101";
			tmp(20,10) := "00010100";
			tmp(20,11) := "01110110";
			tmp(20,12) := "11100011";
			tmp(20,13) := "11101111";
			tmp(20,14) := "11110110";
			tmp(20,15) := "11110111";
			tmp(20,16) := "11101010";
			tmp(20,17) := "11001001";
			tmp(20,18) := "01000000";
			tmp(20,19) := "00010100";
			tmp(20,20) := "01001110";
			tmp(20,21) := "10001110";
			tmp(20,22) := "10011001";
			tmp(20,23) := "10001100";
			tmp(20,24) := "10010101";
			tmp(20,25) := "10011010";
			tmp(20,26) := "10010110";
			tmp(20,27) := "10001011";
			tmp(20,28) := "10001000";
			tmp(20,29) := "10000101";
			tmp(20,30) := "10000011";
			tmp(20,31) := "10000001";
			tmp(20,32) := "01111111";
			tmp(20,33) := "01111100";
			tmp(20,34) := "01111010";
			tmp(20,35) := "01110111";
			tmp(20,36) := "01110100";
			tmp(20,37) := "01110001";
			tmp(20,38) := "01101110";
			tmp(20,39) := "01101011";
			tmp(20,40) := "01101000";
			tmp(21,1) := "10000100";
			tmp(21,2) := "01111110";
			tmp(21,3) := "01111111";
			tmp(21,4) := "01110000";
			tmp(21,5) := "10000000";
			tmp(21,6) := "10000001";
			tmp(21,7) := "01111111";
			tmp(21,8) := "01111101";
			tmp(21,9) := "10000011";
			tmp(21,10) := "10001001";
			tmp(21,11) := "10000000";
			tmp(21,12) := "01111110";
			tmp(21,13) := "01111110";
			tmp(21,14) := "01111001";
			tmp(21,15) := "01111000";
			tmp(21,16) := "01111000";
			tmp(21,17) := "01110110";
			tmp(21,18) := "01111101";
			tmp(21,19) := "10001000";
			tmp(21,20) := "10010001";
			tmp(21,21) := "10011001";
			tmp(21,22) := "10011111";
			tmp(21,23) := "10010110";
			tmp(21,24) := "10001110";
			tmp(21,25) := "10010001";
			tmp(21,26) := "10010010";
			tmp(21,27) := "10001010";
			tmp(21,28) := "10000111";
			tmp(21,29) := "10000100";
			tmp(21,30) := "10000010";
			tmp(21,31) := "10000001";
			tmp(21,32) := "01111110";
			tmp(21,33) := "01111011";
			tmp(21,34) := "01111001";
			tmp(21,35) := "01110110";
			tmp(21,36) := "01110011";
			tmp(21,37) := "01110000";
			tmp(21,38) := "01101101";
			tmp(21,39) := "01101010";
			tmp(21,40) := "01100111";
			tmp(22,1) := "11010000";
			tmp(22,2) := "01011001";
			tmp(22,3) := "00010001";
			tmp(22,4) := "00000000";
			tmp(22,5) := "00011000";
			tmp(22,6) := "01101110";
			tmp(22,7) := "11100010";
			tmp(22,8) := "11110110";
			tmp(22,9) := "11110011";
			tmp(22,10) := "11101110";
			tmp(22,11) := "10010100";
			tmp(22,12) := "00011011";
			tmp(22,13) := "00001010";
			tmp(22,14) := "00000101";
			tmp(22,15) := "00000101";
			tmp(22,16) := "00001001";
			tmp(22,17) := "00101000";
			tmp(22,18) := "10111111";
			tmp(22,19) := "11110001";
			tmp(22,20) := "11001001";
			tmp(22,21) := "10010111";
			tmp(22,22) := "10010100";
			tmp(22,23) := "10011100";
			tmp(22,24) := "10010101";
			tmp(22,25) := "10010101";
			tmp(22,26) := "10001110";
			tmp(22,27) := "10001000";
			tmp(22,28) := "10000110";
			tmp(22,29) := "10000011";
			tmp(22,30) := "10000001";
			tmp(22,31) := "01111111";
			tmp(22,32) := "01111101";
			tmp(22,33) := "01111010";
			tmp(22,34) := "01110111";
			tmp(22,35) := "01110101";
			tmp(22,36) := "01110011";
			tmp(22,37) := "01101111";
			tmp(22,38) := "01101100";
			tmp(22,39) := "01101010";
			tmp(22,40) := "01100111";
			tmp(23,1) := "11010110";
			tmp(23,2) := "01010100";
			tmp(23,3) := "00001010";
			tmp(23,4) := "00000000";
			tmp(23,5) := "00000110";
			tmp(23,6) := "01011110";
			tmp(23,7) := "11111100";
			tmp(23,8) := "11111111";
			tmp(23,9) := "11111100";
			tmp(23,10) := "11110001";
			tmp(23,11) := "10010110";
			tmp(23,12) := "00000111";
			tmp(23,13) := "00000010";
			tmp(23,14) := "00001001";
			tmp(23,15) := "00001011";
			tmp(23,16) := "00000001";
			tmp(23,17) := "00010110";
			tmp(23,18) := "11001011";
			tmp(23,19) := "11111111";
			tmp(23,20) := "11011100";
			tmp(23,21) := "10010110";
			tmp(23,22) := "10001100";
			tmp(23,23) := "10011000";
			tmp(23,24) := "10010110";
			tmp(23,25) := "10011011";
			tmp(23,26) := "10001101";
			tmp(23,27) := "10000111";
			tmp(23,28) := "10000101";
			tmp(23,29) := "10000010";
			tmp(23,30) := "10000000";
			tmp(23,31) := "01111110";
			tmp(23,32) := "01111100";
			tmp(23,33) := "01111001";
			tmp(23,34) := "01111000";
			tmp(23,35) := "01110101";
			tmp(23,36) := "01110010";
			tmp(23,37) := "01101110";
			tmp(23,38) := "01101011";
			tmp(23,39) := "01101001";
			tmp(23,40) := "01100110";
			tmp(24,1) := "11100010";
			tmp(24,2) := "01001001";
			tmp(24,3) := "00000000";
			tmp(24,4) := "00000000";
			tmp(24,5) := "00000101";
			tmp(24,6) := "01001001";
			tmp(24,7) := "11101110";
			tmp(24,8) := "11111110";
			tmp(24,9) := "11111011";
			tmp(24,10) := "11111110";
			tmp(24,11) := "10011010";
			tmp(24,12) := "00011001";
			tmp(24,13) := "00000101";
			tmp(24,14) := "00000000";
			tmp(24,15) := "00000000";
			tmp(24,16) := "00000001";
			tmp(24,17) := "00011101";
			tmp(24,18) := "11000011";
			tmp(24,19) := "11111001";
			tmp(24,20) := "11100111";
			tmp(24,21) := "10101010";
			tmp(24,22) := "10010101";
			tmp(24,23) := "10010101";
			tmp(24,24) := "10010000";
			tmp(24,25) := "10011000";
			tmp(24,26) := "10000111";
			tmp(24,27) := "10000110";
			tmp(24,28) := "10000100";
			tmp(24,29) := "10000001";
			tmp(24,30) := "01111111";
			tmp(24,31) := "01111101";
			tmp(24,32) := "01111011";
			tmp(24,33) := "01111000";
			tmp(24,34) := "01110110";
			tmp(24,35) := "01110100";
			tmp(24,36) := "01110010";
			tmp(24,37) := "01101110";
			tmp(24,38) := "01101011";
			tmp(24,39) := "01101001";
			tmp(24,40) := "01100110";
			tmp(25,1) := "11101000";
			tmp(25,2) := "01010111";
			tmp(25,3) := "00000010";
			tmp(25,4) := "00000000";
			tmp(25,5) := "00000111";
			tmp(25,6) := "01001100";
			tmp(25,7) := "11110010";
			tmp(25,8) := "11111101";
			tmp(25,9) := "11111110";
			tmp(25,10) := "11111110";
			tmp(25,11) := "10100011";
			tmp(25,12) := "00010111";
			tmp(25,13) := "00000001";
			tmp(25,14) := "00000000";
			tmp(25,15) := "00000000";
			tmp(25,16) := "00000000";
			tmp(25,17) := "00011001";
			tmp(25,18) := "10110110";
			tmp(25,19) := "11111111";
			tmp(25,20) := "11101110";
			tmp(25,21) := "10111011";
			tmp(25,22) := "10010111";
			tmp(25,23) := "10011000";
			tmp(25,24) := "10001110";
			tmp(25,25) := "10000101";
			tmp(25,26) := "10010011";
			tmp(25,27) := "10000011";
			tmp(25,28) := "10000001";
			tmp(25,29) := "01111111";
			tmp(25,30) := "01111101";
			tmp(25,31) := "01111100";
			tmp(25,32) := "01111010";
			tmp(25,33) := "01110111";
			tmp(25,34) := "01110101";
			tmp(25,35) := "01110001";
			tmp(25,36) := "01101110";
			tmp(25,37) := "01101010";
			tmp(25,38) := "01101000";
			tmp(25,39) := "01100111";
			tmp(25,40) := "01100101";
			tmp(26,1) := "11101000";
			tmp(26,2) := "01010111";
			tmp(26,3) := "00000010";
			tmp(26,4) := "00000000";
			tmp(26,5) := "00000110";
			tmp(26,6) := "01001010";
			tmp(26,7) := "11110001";
			tmp(26,8) := "11111101";
			tmp(26,9) := "11111110";
			tmp(26,10) := "11111110";
			tmp(26,11) := "10100101";
			tmp(26,12) := "00011000";
			tmp(26,13) := "00000001";
			tmp(26,14) := "00000000";
			tmp(26,15) := "00000000";
			tmp(26,16) := "00000000";
			tmp(26,17) := "00011000";
			tmp(26,18) := "10110100";
			tmp(26,19) := "11111111";
			tmp(26,20) := "11110111";
			tmp(26,21) := "11001011";
			tmp(26,22) := "10011100";
			tmp(26,23) := "10010010";
			tmp(26,24) := "10010100";
			tmp(26,25) := "10001110";
			tmp(26,26) := "10001010";
			tmp(26,27) := "10000010";
			tmp(26,28) := "10000000";
			tmp(26,29) := "01111110";
			tmp(26,30) := "01111100";
			tmp(26,31) := "01111011";
			tmp(26,32) := "01111001";
			tmp(26,33) := "01110110";
			tmp(26,34) := "01110100";
			tmp(26,35) := "01110000";
			tmp(26,36) := "01101101";
			tmp(26,37) := "01101001";
			tmp(26,38) := "01101000";
			tmp(26,39) := "01100110";
			tmp(26,40) := "01100101";
			tmp(27,1) := "11101001";
			tmp(27,2) := "01011001";
			tmp(27,3) := "00000010";
			tmp(27,4) := "00000000";
			tmp(27,5) := "00000101";
			tmp(27,6) := "01000111";
			tmp(27,7) := "11101111";
			tmp(27,8) := "11111101";
			tmp(27,9) := "11111111";
			tmp(27,10) := "11111101";
			tmp(27,11) := "10101000";
			tmp(27,12) := "00011001";
			tmp(27,13) := "00000001";
			tmp(27,14) := "00000000";
			tmp(27,15) := "00000000";
			tmp(27,16) := "00000000";
			tmp(27,17) := "00010101";
			tmp(27,18) := "10110000";
			tmp(27,19) := "11111101";
			tmp(27,20) := "11111111";
			tmp(27,21) := "11100011";
			tmp(27,22) := "10101011";
			tmp(27,23) := "10001101";
			tmp(27,24) := "10010101";
			tmp(27,25) := "10010101";
			tmp(27,26) := "10000011";
			tmp(27,27) := "10000001";
			tmp(27,28) := "01111111";
			tmp(27,29) := "01111011";
			tmp(27,30) := "01111010";
			tmp(27,31) := "01111001";
			tmp(27,32) := "01110111";
			tmp(27,33) := "01110100";
			tmp(27,34) := "01110010";
			tmp(27,35) := "01101111";
			tmp(27,36) := "01101100";
			tmp(27,37) := "01101000";
			tmp(27,38) := "01100110";
			tmp(27,39) := "01100100";
			tmp(27,40) := "01100100";
			tmp(28,1) := "11101100";
			tmp(28,2) := "01011100";
			tmp(28,3) := "00000011";
			tmp(28,4) := "00000000";
			tmp(28,5) := "00000011";
			tmp(28,6) := "01000011";
			tmp(28,7) := "11101100";
			tmp(28,8) := "11111101";
			tmp(28,9) := "11111111";
			tmp(28,10) := "11111100";
			tmp(28,11) := "10101100";
			tmp(28,12) := "00011011";
			tmp(28,13) := "00000001";
			tmp(28,14) := "00000000";
			tmp(28,15) := "00000001";
			tmp(28,16) := "00000000";
			tmp(28,17) := "00010010";
			tmp(28,18) := "10101010";
			tmp(28,19) := "11111101";
			tmp(28,20) := "11111110";
			tmp(28,21) := "11110111";
			tmp(28,22) := "11000100";
			tmp(28,23) := "10010100";
			tmp(28,24) := "10001111";
			tmp(28,25) := "10010011";
			tmp(28,26) := "10000100";
			tmp(28,27) := "10000000";
			tmp(28,28) := "01111101";
			tmp(28,29) := "01111010";
			tmp(28,30) := "01110111";
			tmp(28,31) := "01110110";
			tmp(28,32) := "01110100";
			tmp(28,33) := "01110010";
			tmp(28,34) := "01110000";
			tmp(28,35) := "01101100";
			tmp(28,36) := "01101010";
			tmp(28,37) := "01100110";
			tmp(28,38) := "01100100";
			tmp(28,39) := "01100011";
			tmp(28,40) := "01100010";
			tmp(29,1) := "11101110";
			tmp(29,2) := "01100001";
			tmp(29,3) := "00000100";
			tmp(29,4) := "00000000";
			tmp(29,5) := "00000001";
			tmp(29,6) := "00111111";
			tmp(29,7) := "11101000";
			tmp(29,8) := "11111100";
			tmp(29,9) := "11111111";
			tmp(29,10) := "11111011";
			tmp(29,11) := "10101111";
			tmp(29,12) := "00011101";
			tmp(29,13) := "00000010";
			tmp(29,14) := "00000000";
			tmp(29,15) := "00000001";
			tmp(29,16) := "00000000";
			tmp(29,17) := "00001111";
			tmp(29,18) := "10100100";
			tmp(29,19) := "11111100";
			tmp(29,20) := "11111111";
			tmp(29,21) := "11111111";
			tmp(29,22) := "11100000";
			tmp(29,23) := "10101010";
			tmp(29,24) := "10001011";
			tmp(29,25) := "10001010";
			tmp(29,26) := "10001100";
			tmp(29,27) := "01111111";
			tmp(29,28) := "01111100";
			tmp(29,29) := "01110111";
			tmp(29,30) := "01110100";
			tmp(29,31) := "01110011";
			tmp(29,32) := "01110001";
			tmp(29,33) := "01101111";
			tmp(29,34) := "01101101";
			tmp(29,35) := "01101010";
			tmp(29,36) := "01101000";
			tmp(29,37) := "01100100";
			tmp(29,38) := "01100010";
			tmp(29,39) := "01100010";
			tmp(29,40) := "01100001";
			tmp(30,1) := "11110001";
			tmp(30,2) := "01100100";
			tmp(30,3) := "00000101";
			tmp(30,4) := "00000000";
			tmp(30,5) := "00000000";
			tmp(30,6) := "00111011";
			tmp(30,7) := "11100101";
			tmp(30,8) := "11111100";
			tmp(30,9) := "11111111";
			tmp(30,10) := "11111011";
			tmp(30,11) := "10110011";
			tmp(30,12) := "00011110";
			tmp(30,13) := "00000010";
			tmp(30,14) := "00000000";
			tmp(30,15) := "00000010";
			tmp(30,16) := "00000000";
			tmp(30,17) := "00001100";
			tmp(30,18) := "10011111";
			tmp(30,19) := "11111011";
			tmp(30,20) := "11111100";
			tmp(30,21) := "11111111";
			tmp(30,22) := "11110101";
			tmp(30,23) := "11001000";
			tmp(30,24) := "10010111";
			tmp(30,25) := "10000110";
			tmp(30,26) := "10001111";
			tmp(30,27) := "01111110";
			tmp(30,28) := "01111010";
			tmp(30,29) := "01110101";
			tmp(30,30) := "01110001";
			tmp(30,31) := "01110000";
			tmp(30,32) := "01101110";
			tmp(30,33) := "01101101";
			tmp(30,34) := "01101011";
			tmp(30,35) := "01101000";
			tmp(30,36) := "01100110";
			tmp(30,37) := "01100010";
			tmp(30,38) := "01100001";
			tmp(30,39) := "01100000";
			tmp(30,40) := "01100000";
			tmp(31,1) := "11110010";
			tmp(31,2) := "01100110";
			tmp(31,3) := "00000101";
			tmp(31,4) := "00000000";
			tmp(31,5) := "00000000";
			tmp(31,6) := "00111000";
			tmp(31,7) := "11100011";
			tmp(31,8) := "11111011";
			tmp(31,9) := "11111111";
			tmp(31,10) := "11111010";
			tmp(31,11) := "10110101";
			tmp(31,12) := "00100000";
			tmp(31,13) := "00000010";
			tmp(31,14) := "00000000";
			tmp(31,15) := "00000010";
			tmp(31,16) := "00000000";
			tmp(31,17) := "00001010";
			tmp(31,18) := "10011011";
			tmp(31,19) := "11111010";
			tmp(31,20) := "11111111";
			tmp(31,21) := "11111110";
			tmp(31,22) := "11111101";
			tmp(31,23) := "11100110";
			tmp(31,24) := "10110001";
			tmp(31,25) := "10001010";
			tmp(31,26) := "10001100";
			tmp(31,27) := "01111101";
			tmp(31,28) := "01111001";
			tmp(31,29) := "01110011";
			tmp(31,30) := "01101111";
			tmp(31,31) := "01101101";
			tmp(31,32) := "01101100";
			tmp(31,33) := "01101011";
			tmp(31,34) := "01101010";
			tmp(31,35) := "01100111";
			tmp(31,36) := "01100100";
			tmp(31,37) := "01100001";
			tmp(31,38) := "01011111";
			tmp(31,39) := "01011111";
			tmp(31,40) := "01011110";
			tmp(32,1) := "11110010";
			tmp(32,2) := "01100110";
			tmp(32,3) := "00000101";
			tmp(32,4) := "00000000";
			tmp(32,5) := "00000001";
			tmp(32,6) := "00110110";
			tmp(32,7) := "11100001";
			tmp(32,8) := "11111011";
			tmp(32,9) := "11111111";
			tmp(32,10) := "11111010";
			tmp(32,11) := "10110111";
			tmp(32,12) := "00100001";
			tmp(32,13) := "00000010";
			tmp(32,14) := "00000000";
			tmp(32,15) := "00000010";
			tmp(32,16) := "00000000";
			tmp(32,17) := "00001000";
			tmp(32,18) := "10011000";
			tmp(32,19) := "11111001";
			tmp(32,20) := "11111111";
			tmp(32,21) := "11111110";
			tmp(32,22) := "11111101";
			tmp(32,23) := "11111000";
			tmp(32,24) := "11000110";
			tmp(32,25) := "10010000";
			tmp(32,26) := "10000110";
			tmp(32,27) := "01111100";
			tmp(32,28) := "01111000";
			tmp(32,29) := "01110010";
			tmp(32,30) := "01101110";
			tmp(32,31) := "01101100";
			tmp(32,32) := "01101011";
			tmp(32,33) := "01101010";
			tmp(32,34) := "01101001";
			tmp(32,35) := "01100110";
			tmp(32,36) := "01100011";
			tmp(32,37) := "01100000";
			tmp(32,38) := "01011111";
			tmp(32,39) := "01011111";
			tmp(32,40) := "01011110";
			tmp(33,1) := "11101111";
			tmp(33,2) := "01111000";
			tmp(33,3) := "00001001";
			tmp(33,4) := "00000000";
			tmp(33,5) := "00001011";
			tmp(33,6) := "00111111";
			tmp(33,7) := "11010111";
			tmp(33,8) := "11111101";
			tmp(33,9) := "11111111";
			tmp(33,10) := "11111100";
			tmp(33,11) := "10111011";
			tmp(33,12) := "00101111";
			tmp(33,13) := "00000000";
			tmp(33,14) := "00001001";
			tmp(33,15) := "00000000";
			tmp(33,16) := "00000001";
			tmp(33,17) := "00010110";
			tmp(33,18) := "10011001";
			tmp(33,19) := "11111101";
			tmp(33,20) := "11111111";
			tmp(33,21) := "11111110";
			tmp(33,22) := "11111000";
			tmp(33,23) := "11111111";
			tmp(33,24) := "11101111";
			tmp(33,25) := "10110101";
			tmp(33,26) := "10010100";
			tmp(33,27) := "10000100";
			tmp(33,28) := "01110111";
			tmp(33,29) := "01101101";
			tmp(33,30) := "01101101";
			tmp(33,31) := "01101011";
			tmp(33,32) := "01100011";
			tmp(33,33) := "01100001";
			tmp(33,34) := "01100110";
			tmp(33,35) := "01100000";
			tmp(33,36) := "01100000";
			tmp(33,37) := "01011111";
			tmp(33,38) := "01011110";
			tmp(33,39) := "01011101";
			tmp(33,40) := "01011011";
			tmp(34,1) := "11111011";
			tmp(34,2) := "01100010";
			tmp(34,3) := "00001100";
			tmp(34,4) := "00000000";
			tmp(34,5) := "00000000";
			tmp(34,6) := "00100111";
			tmp(34,7) := "11011010";
			tmp(34,8) := "11111111";
			tmp(34,9) := "11111011";
			tmp(34,10) := "11111010";
			tmp(34,11) := "11000010";
			tmp(34,12) := "00110000";
			tmp(34,13) := "00000000";
			tmp(34,14) := "00001101";
			tmp(34,15) := "00000000";
			tmp(34,16) := "00000000";
			tmp(34,17) := "00000011";
			tmp(34,18) := "01111011";
			tmp(34,19) := "11111111";
			tmp(34,20) := "11111100";
			tmp(34,21) := "11111100";
			tmp(34,22) := "11110111";
			tmp(34,23) := "11111111";
			tmp(34,24) := "11111011";
			tmp(34,25) := "11001010";
			tmp(34,26) := "10011010";
			tmp(34,27) := "10000001";
			tmp(34,28) := "01110110";
			tmp(34,29) := "01101101";
			tmp(34,30) := "01101011";
			tmp(34,31) := "01101011";
			tmp(34,32) := "01100110";
			tmp(34,33) := "01011111";
			tmp(34,34) := "01011011";
			tmp(34,35) := "01011110";
			tmp(34,36) := "01011110";
			tmp(34,37) := "01011101";
			tmp(34,38) := "01011100";
			tmp(34,39) := "01011010";
			tmp(34,40) := "01011010";
			tmp(35,1) := "11010001";
			tmp(35,2) := "01110110";
			tmp(35,3) := "00000100";
			tmp(35,4) := "00001100";
			tmp(35,5) := "00000000";
			tmp(35,6) := "00101110";
			tmp(35,7) := "11011000";
			tmp(35,8) := "11111111";
			tmp(35,9) := "11110101";
			tmp(35,10) := "11111111";
			tmp(35,11) := "11000101";
			tmp(35,12) := "00100000";
			tmp(35,13) := "00000000";
			tmp(35,14) := "00000011";
			tmp(35,15) := "00000000";
			tmp(35,16) := "00001110";
			tmp(35,17) := "00001101";
			tmp(35,18) := "10000110";
			tmp(35,19) := "11111111";
			tmp(35,20) := "11111000";
			tmp(35,21) := "11111101";
			tmp(35,22) := "11111100";
			tmp(35,23) := "11111101";
			tmp(35,24) := "11111111";
			tmp(35,25) := "11011001";
			tmp(35,26) := "10000110";
			tmp(35,27) := "01110101";
			tmp(35,28) := "01110101";
			tmp(35,29) := "01101111";
			tmp(35,30) := "01100100";
			tmp(35,31) := "01011101";
			tmp(35,32) := "01011011";
			tmp(35,33) := "01011110";
			tmp(35,34) := "01011111";
			tmp(35,35) := "01011011";
			tmp(35,36) := "01011011";
			tmp(35,37) := "01011010";
			tmp(35,38) := "01011001";
			tmp(35,39) := "01011000";
			tmp(35,40) := "01010111";
			tmp(36,1) := "01001000";
			tmp(36,2) := "01101100";
			tmp(36,3) := "01011001";
			tmp(36,4) := "01000001";
			tmp(36,5) := "00010100";
			tmp(36,6) := "00111111";
			tmp(36,7) := "11001111";
			tmp(36,8) := "11111111";
			tmp(36,9) := "11110111";
			tmp(36,10) := "11111100";
			tmp(36,11) := "11000101";
			tmp(36,12) := "00101001";
			tmp(36,13) := "00000110";
			tmp(36,14) := "00001010";
			tmp(36,15) := "00000000";
			tmp(36,16) := "00000000";
			tmp(36,17) := "00000000";
			tmp(36,18) := "10001110";
			tmp(36,19) := "11111011";
			tmp(36,20) := "11110111";
			tmp(36,21) := "11111111";
			tmp(36,22) := "11111111";
			tmp(36,23) := "11111100";
			tmp(36,24) := "11111111";
			tmp(36,25) := "11010111";
			tmp(36,26) := "01011111";
			tmp(36,27) := "01000110";
			tmp(36,28) := "01011111";
			tmp(36,29) := "01110000";
			tmp(36,30) := "01101001";
			tmp(36,31) := "01011011";
			tmp(36,32) := "01010111";
			tmp(36,33) := "01011010";
			tmp(36,34) := "01011101";
			tmp(36,35) := "01011000";
			tmp(36,36) := "01011000";
			tmp(36,37) := "01010111";
			tmp(36,38) := "01010110";
			tmp(36,39) := "01010101";
			tmp(36,40) := "01010101";
			tmp(37,1) := "00001100";
			tmp(37,2) := "01110101";
			tmp(37,3) := "11100110";
			tmp(37,4) := "11000111";
			tmp(37,5) := "10011111";
			tmp(37,6) := "10011010";
			tmp(37,7) := "10101001";
			tmp(37,8) := "11001001";
			tmp(37,9) := "11100001";
			tmp(37,10) := "11111010";
			tmp(37,11) := "11001011";
			tmp(37,12) := "00110011";
			tmp(37,13) := "00000000";
			tmp(37,14) := "00000101";
			tmp(37,15) := "00000110";
			tmp(37,16) := "00001100";
			tmp(37,17) := "00000000";
			tmp(37,18) := "01111101";
			tmp(37,19) := "11111100";
			tmp(37,20) := "11111011";
			tmp(37,21) := "11111111";
			tmp(37,22) := "11111111";
			tmp(37,23) := "11111000";
			tmp(37,24) := "11111110";
			tmp(37,25) := "11010111";
			tmp(37,26) := "01001010";
			tmp(37,27) := "00001100";
			tmp(37,28) := "00110000";
			tmp(37,29) := "01010101";
			tmp(37,30) := "01100101";
			tmp(37,31) := "01100110";
			tmp(37,32) := "01100001";
			tmp(37,33) := "01011001";
			tmp(37,34) := "01001111";
			tmp(37,35) := "01010101";
			tmp(37,36) := "01010101";
			tmp(37,37) := "01010100";
			tmp(37,38) := "01010100";
			tmp(37,39) := "01010011";
			tmp(37,40) := "01010010";
			tmp(38,1) := "00000110";
			tmp(38,2) := "01111010";
			tmp(38,3) := "11110001";
			tmp(38,4) := "11111110";
			tmp(38,5) := "11111111";
			tmp(38,6) := "11010101";
			tmp(38,7) := "01001010";
			tmp(38,8) := "00101001";
			tmp(38,9) := "01010110";
			tmp(38,10) := "10000110";
			tmp(38,11) := "10010010";
			tmp(38,12) := "00111110";
			tmp(38,13) := "00000011";
			tmp(38,14) := "00000000";
			tmp(38,15) := "00000000";
			tmp(38,16) := "00000100";
			tmp(38,17) := "00000000";
			tmp(38,18) := "01101110";
			tmp(38,19) := "11111101";
			tmp(38,20) := "11111111";
			tmp(38,21) := "11111101";
			tmp(38,22) := "11111111";
			tmp(38,23) := "11110101";
			tmp(38,24) := "11111111";
			tmp(38,25) := "11100001";
			tmp(38,26) := "01010011";
			tmp(38,27) := "00000000";
			tmp(38,28) := "00001011";
			tmp(38,29) := "00011110";
			tmp(38,30) := "00110101";
			tmp(38,31) := "01001101";
			tmp(38,32) := "01011011";
			tmp(38,33) := "01011010";
			tmp(38,34) := "01010010";
			tmp(38,35) := "01010000";
			tmp(38,36) := "01010000";
			tmp(38,37) := "01010000";
			tmp(38,38) := "01001111";
			tmp(38,39) := "01001111";
			tmp(38,40) := "01001101";
			tmp(39,1) := "00001111";
			tmp(39,2) := "01111100";
			tmp(39,3) := "11110001";
			tmp(39,4) := "11111011";
			tmp(39,5) := "11111111";
			tmp(39,6) := "11011110";
			tmp(39,7) := "00110101";
			tmp(39,8) := "00000000";
			tmp(39,9) := "00000000";
			tmp(39,10) := "00001001";
			tmp(39,11) := "00110100";
			tmp(39,12) := "10000000";
			tmp(39,13) := "10000000";
			tmp(39,14) := "01010101";
			tmp(39,15) := "00011110";
			tmp(39,16) := "00000010";
			tmp(39,17) := "00001011";
			tmp(39,18) := "01110100";
			tmp(39,19) := "11110101";
			tmp(39,20) := "11111111";
			tmp(39,21) := "11111010";
			tmp(39,22) := "11111111";
			tmp(39,23) := "11111000";
			tmp(39,24) := "11111111";
			tmp(39,25) := "11100101";
			tmp(39,26) := "01011101";
			tmp(39,27) := "00001011";
			tmp(39,28) := "00000000";
			tmp(39,29) := "00000000";
			tmp(39,30) := "00000111";
			tmp(39,31) := "00011111";
			tmp(39,32) := "00110110";
			tmp(39,33) := "01001001";
			tmp(39,34) := "01010100";
			tmp(39,35) := "01001011";
			tmp(39,36) := "01001011";
			tmp(39,37) := "01001010";
			tmp(39,38) := "01001010";
			tmp(39,39) := "01001010";
			tmp(39,40) := "01001001";
			tmp(40,1) := "00010001";
			tmp(40,2) := "01101110";
			tmp(40,3) := "11110110";
			tmp(40,4) := "11111010";
			tmp(40,5) := "11111110";
			tmp(40,6) := "11011011";
			tmp(40,7) := "00111001";
			tmp(40,8) := "00000101";
			tmp(40,9) := "00000000";
			tmp(40,10) := "00000001";
			tmp(40,11) := "00100111";
			tmp(40,12) := "11001011";
			tmp(40,13) := "11110101";
			tmp(40,14) := "11100011";
			tmp(40,15) := "11000110";
			tmp(40,16) := "10011011";
			tmp(40,17) := "01101101";
			tmp(40,18) := "10001010";
			tmp(40,19) := "11101000";
			tmp(40,20) := "11111110";
			tmp(40,21) := "11111001";
			tmp(40,22) := "11111111";
			tmp(40,23) := "11111111";
			tmp(40,24) := "11111111";
			tmp(40,25) := "11100000";
			tmp(40,26) := "01011011";
			tmp(40,27) := "00000100";
			tmp(40,28) := "00000000";
			tmp(40,29) := "00000000";
			tmp(40,30) := "00000011";
			tmp(40,31) := "00001010";
			tmp(40,32) := "00010100";
			tmp(40,33) := "00101010";
			tmp(40,34) := "01000001";
			tmp(40,35) := "01000110";
			tmp(40,36) := "01000110";
			tmp(40,37) := "01000110";
			tmp(40,38) := "01000110";
			tmp(40,39) := "01000110";
			tmp(40,40) := "01000101";

		return tmp;
	end init_rom;
	
	-- Declare the ROM signal and specify a default value.	Quartus II
	-- will create a memory initialization file (.mif) based on the 
	-- default value.
	signal rom : memory_t := init_rom;
begin
	process(clk)
	variable t : matrix_in;
	begin
		for i in addr_i to (addr_i + elin-1) loop
			for j in addr_j to (addr_j + ecol-1) loop
				t(i-addr_i, j-addr_j) := rom(addr_i+(i-addr_i), addr_j+(j-addr_j));
			end loop;
		end loop;
		if(rising_edge(clk)) then
			q <= t;
		end if;
	end process;
		
end rtl;
