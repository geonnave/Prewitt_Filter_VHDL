library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.mem_size.all;
use work.matrix_types.all;

entity MemImgROM is
	port
	(
		addr_i	:	in	natural		range 0 to lin-1;
		addr_j	:	in	natural		range 0 to col-1;
		clk		:	in std_logic;
		q		:	out matrix_in
	);
end entity;


architecture rtl of MemImgROM is

	-- Build a 2-D array type for the RoM
	subtype pixel is std_logic_vector(7 downto 0);
	type memory_t is array(0 to lin, 0 to col) of pixel;
		
	function init_rom
		return memory_t is
		variable tmp : memory_t;
		begin
			tmp(0,0) := "00000000";
			tmp(81,0) := "00000000";
			tmp(0,1) := "00000000";
			tmp(81,1) := "00000000";
			tmp(0,2) := "00000000";
			tmp(81,2) := "00000000";
			tmp(0,3) := "00000000";
			tmp(81,3) := "00000000";
			tmp(0,4) := "00000000";
			tmp(81,4) := "00000000";
			tmp(0,5) := "00000000";
			tmp(81,5) := "00000000";
			tmp(0,6) := "00000000";
			tmp(81,6) := "00000000";
			tmp(0,7) := "00000000";
			tmp(81,7) := "00000000";
			tmp(0,8) := "00000000";
			tmp(81,8) := "00000000";
			tmp(0,9) := "00000000";
			tmp(81,9) := "00000000";
			tmp(0,10) := "00000000";
			tmp(81,10) := "00000000";
			tmp(0,11) := "00000000";
			tmp(81,11) := "00000000";
			tmp(0,12) := "00000000";
			tmp(81,12) := "00000000";
			tmp(0,13) := "00000000";
			tmp(81,13) := "00000000";
			tmp(0,14) := "00000000";
			tmp(81,14) := "00000000";
			tmp(0,15) := "00000000";
			tmp(81,15) := "00000000";
			tmp(0,16) := "00000000";
			tmp(81,16) := "00000000";
			tmp(0,17) := "00000000";
			tmp(81,17) := "00000000";
			tmp(0,18) := "00000000";
			tmp(81,18) := "00000000";
			tmp(0,19) := "00000000";
			tmp(81,19) := "00000000";
			tmp(0,20) := "00000000";
			tmp(81,20) := "00000000";
			tmp(0,21) := "00000000";
			tmp(81,21) := "00000000";
			tmp(0,22) := "00000000";
			tmp(81,22) := "00000000";
			tmp(0,23) := "00000000";
			tmp(81,23) := "00000000";
			tmp(0,24) := "00000000";
			tmp(81,24) := "00000000";
			tmp(0,25) := "00000000";
			tmp(81,25) := "00000000";
			tmp(0,26) := "00000000";
			tmp(81,26) := "00000000";
			tmp(0,27) := "00000000";
			tmp(81,27) := "00000000";
			tmp(0,28) := "00000000";
			tmp(81,28) := "00000000";
			tmp(0,29) := "00000000";
			tmp(81,29) := "00000000";
			tmp(0,30) := "00000000";
			tmp(81,30) := "00000000";
			tmp(0,31) := "00000000";
			tmp(81,31) := "00000000";
			tmp(0,32) := "00000000";
			tmp(81,32) := "00000000";
			tmp(0,33) := "00000000";
			tmp(81,33) := "00000000";
			tmp(0,34) := "00000000";
			tmp(81,34) := "00000000";
			tmp(0,35) := "00000000";
			tmp(81,35) := "00000000";
			tmp(0,36) := "00000000";
			tmp(81,36) := "00000000";
			tmp(0,37) := "00000000";
			tmp(81,37) := "00000000";
			tmp(0,38) := "00000000";
			tmp(81,38) := "00000000";
			tmp(0,39) := "00000000";
			tmp(81,39) := "00000000";
			tmp(0,40) := "00000000";
			tmp(81,40) := "00000000";
			tmp(0,41) := "00000000";
			tmp(81,41) := "00000000";
			tmp(0,42) := "00000000";
			tmp(81,42) := "00000000";
			tmp(0,43) := "00000000";
			tmp(81,43) := "00000000";
			tmp(0,44) := "00000000";
			tmp(81,44) := "00000000";
			tmp(0,45) := "00000000";
			tmp(81,45) := "00000000";
			tmp(0,46) := "00000000";
			tmp(81,46) := "00000000";
			tmp(0,47) := "00000000";
			tmp(81,47) := "00000000";
			tmp(0,48) := "00000000";
			tmp(81,48) := "00000000";
			tmp(0,49) := "00000000";
			tmp(81,49) := "00000000";
			tmp(0,50) := "00000000";
			tmp(81,50) := "00000000";
			tmp(0,51) := "00000000";
			tmp(81,51) := "00000000";
			tmp(0,52) := "00000000";
			tmp(81,52) := "00000000";
			tmp(0,53) := "00000000";
			tmp(81,53) := "00000000";
			tmp(0,54) := "00000000";
			tmp(81,54) := "00000000";
			tmp(0,55) := "00000000";
			tmp(81,55) := "00000000";
			tmp(0,56) := "00000000";
			tmp(81,56) := "00000000";
			tmp(0,57) := "00000000";
			tmp(81,57) := "00000000";
			tmp(0,58) := "00000000";
			tmp(81,58) := "00000000";
			tmp(0,59) := "00000000";
			tmp(81,59) := "00000000";
			tmp(0,60) := "00000000";
			tmp(81,60) := "00000000";
			tmp(0,61) := "00000000";
			tmp(81,61) := "00000000";
			tmp(0,62) := "00000000";
			tmp(81,62) := "00000000";
			tmp(0,63) := "00000000";
			tmp(81,63) := "00000000";
			tmp(0,64) := "00000000";
			tmp(81,64) := "00000000";
			tmp(0,65) := "00000000";
			tmp(81,65) := "00000000";
			tmp(0,66) := "00000000";
			tmp(81,66) := "00000000";
			tmp(0,67) := "00000000";
			tmp(81,67) := "00000000";
			tmp(0,68) := "00000000";
			tmp(81,68) := "00000000";
			tmp(0,69) := "00000000";
			tmp(81,69) := "00000000";
			tmp(0,70) := "00000000";
			tmp(81,70) := "00000000";
			tmp(0,71) := "00000000";
			tmp(81,71) := "00000000";
			tmp(0,72) := "00000000";
			tmp(81,72) := "00000000";
			tmp(0,73) := "00000000";
			tmp(81,73) := "00000000";
			tmp(0,74) := "00000000";
			tmp(81,74) := "00000000";
			tmp(0,75) := "00000000";
			tmp(81,75) := "00000000";
			tmp(0,76) := "00000000";
			tmp(81,76) := "00000000";
			tmp(0,77) := "00000000";
			tmp(81,77) := "00000000";
			tmp(0,78) := "00000000";
			tmp(81,78) := "00000000";
			tmp(0,79) := "00000000";
			tmp(81,79) := "00000000";
			tmp(0,80) := "00000000";
			tmp(81,80) := "00000000";
			tmp(0,81) := "00000000";
			tmp(81,81) := "00000000";
			tmp(0,0) := "00000000";
			tmp(0,81) := "00000000";
			tmp(1,0) := "00000000";
			tmp(1,81) := "00000000";
			tmp(2,0) := "00000000";
			tmp(2,81) := "00000000";
			tmp(3,0) := "00000000";
			tmp(3,81) := "00000000";
			tmp(4,0) := "00000000";
			tmp(4,81) := "00000000";
			tmp(5,0) := "00000000";
			tmp(5,81) := "00000000";
			tmp(6,0) := "00000000";
			tmp(6,81) := "00000000";
			tmp(7,0) := "00000000";
			tmp(7,81) := "00000000";
			tmp(8,0) := "00000000";
			tmp(8,81) := "00000000";
			tmp(9,0) := "00000000";
			tmp(9,81) := "00000000";
			tmp(10,0) := "00000000";
			tmp(10,81) := "00000000";
			tmp(11,0) := "00000000";
			tmp(11,81) := "00000000";
			tmp(12,0) := "00000000";
			tmp(12,81) := "00000000";
			tmp(13,0) := "00000000";
			tmp(13,81) := "00000000";
			tmp(14,0) := "00000000";
			tmp(14,81) := "00000000";
			tmp(15,0) := "00000000";
			tmp(15,81) := "00000000";
			tmp(16,0) := "00000000";
			tmp(16,81) := "00000000";
			tmp(17,0) := "00000000";
			tmp(17,81) := "00000000";
			tmp(18,0) := "00000000";
			tmp(18,81) := "00000000";
			tmp(19,0) := "00000000";
			tmp(19,81) := "00000000";
			tmp(20,0) := "00000000";
			tmp(20,81) := "00000000";
			tmp(21,0) := "00000000";
			tmp(21,81) := "00000000";
			tmp(22,0) := "00000000";
			tmp(22,81) := "00000000";
			tmp(23,0) := "00000000";
			tmp(23,81) := "00000000";
			tmp(24,0) := "00000000";
			tmp(24,81) := "00000000";
			tmp(25,0) := "00000000";
			tmp(25,81) := "00000000";
			tmp(26,0) := "00000000";
			tmp(26,81) := "00000000";
			tmp(27,0) := "00000000";
			tmp(27,81) := "00000000";
			tmp(28,0) := "00000000";
			tmp(28,81) := "00000000";
			tmp(29,0) := "00000000";
			tmp(29,81) := "00000000";
			tmp(30,0) := "00000000";
			tmp(30,81) := "00000000";
			tmp(31,0) := "00000000";
			tmp(31,81) := "00000000";
			tmp(32,0) := "00000000";
			tmp(32,81) := "00000000";
			tmp(33,0) := "00000000";
			tmp(33,81) := "00000000";
			tmp(34,0) := "00000000";
			tmp(34,81) := "00000000";
			tmp(35,0) := "00000000";
			tmp(35,81) := "00000000";
			tmp(36,0) := "00000000";
			tmp(36,81) := "00000000";
			tmp(37,0) := "00000000";
			tmp(37,81) := "00000000";
			tmp(38,0) := "00000000";
			tmp(38,81) := "00000000";
			tmp(39,0) := "00000000";
			tmp(39,81) := "00000000";
			tmp(40,0) := "00000000";
			tmp(40,81) := "00000000";
			tmp(41,0) := "00000000";
			tmp(41,81) := "00000000";
			tmp(42,0) := "00000000";
			tmp(42,81) := "00000000";
			tmp(43,0) := "00000000";
			tmp(43,81) := "00000000";
			tmp(44,0) := "00000000";
			tmp(44,81) := "00000000";
			tmp(45,0) := "00000000";
			tmp(45,81) := "00000000";
			tmp(46,0) := "00000000";
			tmp(46,81) := "00000000";
			tmp(47,0) := "00000000";
			tmp(47,81) := "00000000";
			tmp(48,0) := "00000000";
			tmp(48,81) := "00000000";
			tmp(49,0) := "00000000";
			tmp(49,81) := "00000000";
			tmp(50,0) := "00000000";
			tmp(50,81) := "00000000";
			tmp(51,0) := "00000000";
			tmp(51,81) := "00000000";
			tmp(52,0) := "00000000";
			tmp(52,81) := "00000000";
			tmp(53,0) := "00000000";
			tmp(53,81) := "00000000";
			tmp(54,0) := "00000000";
			tmp(54,81) := "00000000";
			tmp(55,0) := "00000000";
			tmp(55,81) := "00000000";
			tmp(56,0) := "00000000";
			tmp(56,81) := "00000000";
			tmp(57,0) := "00000000";
			tmp(57,81) := "00000000";
			tmp(58,0) := "00000000";
			tmp(58,81) := "00000000";
			tmp(59,0) := "00000000";
			tmp(59,81) := "00000000";
			tmp(60,0) := "00000000";
			tmp(60,81) := "00000000";
			tmp(61,0) := "00000000";
			tmp(61,81) := "00000000";
			tmp(62,0) := "00000000";
			tmp(62,81) := "00000000";
			tmp(63,0) := "00000000";
			tmp(63,81) := "00000000";
			tmp(64,0) := "00000000";
			tmp(64,81) := "00000000";
			tmp(65,0) := "00000000";
			tmp(65,81) := "00000000";
			tmp(66,0) := "00000000";
			tmp(66,81) := "00000000";
			tmp(67,0) := "00000000";
			tmp(67,81) := "00000000";
			tmp(68,0) := "00000000";
			tmp(68,81) := "00000000";
			tmp(69,0) := "00000000";
			tmp(69,81) := "00000000";
			tmp(70,0) := "00000000";
			tmp(70,81) := "00000000";
			tmp(71,0) := "00000000";
			tmp(71,81) := "00000000";
			tmp(72,0) := "00000000";
			tmp(72,81) := "00000000";
			tmp(73,0) := "00000000";
			tmp(73,81) := "00000000";
			tmp(74,0) := "00000000";
			tmp(74,81) := "00000000";
			tmp(75,0) := "00000000";
			tmp(75,81) := "00000000";
			tmp(76,0) := "00000000";
			tmp(76,81) := "00000000";
			tmp(77,0) := "00000000";
			tmp(77,81) := "00000000";
			tmp(78,0) := "00000000";
			tmp(78,81) := "00000000";
			tmp(79,0) := "00000000";
			tmp(79,81) := "00000000";
			tmp(80,0) := "00000000";
			tmp(80,81) := "00000000";
			tmp(81,0) := "00000000";
			tmp(81,81) := "00000000";
			tmp(1,1) := "11111111";
			tmp(1,2) := "11111111";
			tmp(1,3) := "11111111";
			tmp(1,4) := "11111111";
			tmp(1,5) := "11111111";
			tmp(1,6) := "11111111";
			tmp(1,7) := "11111111";
			tmp(1,8) := "11111111";
			tmp(1,9) := "11111111";
			tmp(1,10) := "11111111";
			tmp(1,11) := "11111111";
			tmp(1,12) := "11111111";
			tmp(1,13) := "11111111";
			tmp(1,14) := "11111111";
			tmp(1,15) := "11111111";
			tmp(1,16) := "11111111";
			tmp(1,17) := "11111111";
			tmp(1,18) := "11111111";
			tmp(1,19) := "11111111";
			tmp(1,20) := "11111111";
			tmp(1,21) := "11111111";
			tmp(1,22) := "11111111";
			tmp(1,23) := "11111111";
			tmp(1,24) := "11111111";
			tmp(1,25) := "11111111";
			tmp(1,26) := "11111111";
			tmp(1,27) := "11111111";
			tmp(1,28) := "11111111";
			tmp(1,29) := "11111111";
			tmp(1,30) := "11111111";
			tmp(1,31) := "11111111";
			tmp(1,32) := "11111111";
			tmp(1,33) := "11111111";
			tmp(1,34) := "11111111";
			tmp(1,35) := "11111111";
			tmp(1,36) := "11111111";
			tmp(1,37) := "11111111";
			tmp(1,38) := "11111111";
			tmp(1,39) := "11111111";
			tmp(1,40) := "11111111";
			tmp(1,41) := "11111111";
			tmp(1,42) := "11111111";
			tmp(1,43) := "11111111";
			tmp(1,44) := "11111111";
			tmp(1,45) := "11111111";
			tmp(1,46) := "11111111";
			tmp(1,47) := "11111111";
			tmp(1,48) := "11111111";
			tmp(1,49) := "11111111";
			tmp(1,50) := "11111111";
			tmp(1,51) := "11111111";
			tmp(1,52) := "11111111";
			tmp(1,53) := "11111111";
			tmp(1,54) := "11111111";
			tmp(1,55) := "11111111";
			tmp(1,56) := "11111111";
			tmp(1,57) := "11111111";
			tmp(1,58) := "11111111";
			tmp(1,59) := "11111111";
			tmp(1,60) := "11111111";
			tmp(1,61) := "11111111";
			tmp(1,62) := "11111111";
			tmp(1,63) := "11111111";
			tmp(1,64) := "11111111";
			tmp(1,65) := "11111111";
			tmp(1,66) := "11111111";
			tmp(1,67) := "11111111";
			tmp(1,68) := "11111111";
			tmp(1,69) := "11111111";
			tmp(1,70) := "11111111";
			tmp(1,71) := "11111111";
			tmp(1,72) := "11111111";
			tmp(1,73) := "11111111";
			tmp(1,74) := "11111111";
			tmp(1,75) := "11111111";
			tmp(1,76) := "11111111";
			tmp(1,77) := "11111111";
			tmp(1,78) := "11111111";
			tmp(1,79) := "11111111";
			tmp(1,80) := "11111111";
			tmp(2,1) := "11111111";
			tmp(2,2) := "11111111";
			tmp(2,3) := "11111111";
			tmp(2,4) := "11111111";
			tmp(2,5) := "11111111";
			tmp(2,6) := "11111111";
			tmp(2,7) := "11111111";
			tmp(2,8) := "11111111";
			tmp(2,9) := "11111111";
			tmp(2,10) := "11111111";
			tmp(2,11) := "11111111";
			tmp(2,12) := "11111111";
			tmp(2,13) := "11111111";
			tmp(2,14) := "11111111";
			tmp(2,15) := "11111111";
			tmp(2,16) := "11111111";
			tmp(2,17) := "11111111";
			tmp(2,18) := "11111111";
			tmp(2,19) := "11111111";
			tmp(2,20) := "11111111";
			tmp(2,21) := "11111111";
			tmp(2,22) := "11111111";
			tmp(2,23) := "11111111";
			tmp(2,24) := "11111111";
			tmp(2,25) := "11111111";
			tmp(2,26) := "11111111";
			tmp(2,27) := "11111111";
			tmp(2,28) := "11111111";
			tmp(2,29) := "11111111";
			tmp(2,30) := "11111111";
			tmp(2,31) := "11111111";
			tmp(2,32) := "11111111";
			tmp(2,33) := "11111111";
			tmp(2,34) := "11111111";
			tmp(2,35) := "11111111";
			tmp(2,36) := "11111111";
			tmp(2,37) := "11111111";
			tmp(2,38) := "11111111";
			tmp(2,39) := "11111111";
			tmp(2,40) := "11111111";
			tmp(2,41) := "11111111";
			tmp(2,42) := "11111111";
			tmp(2,43) := "11111111";
			tmp(2,44) := "11111111";
			tmp(2,45) := "11111111";
			tmp(2,46) := "11111111";
			tmp(2,47) := "11111111";
			tmp(2,48) := "11111111";
			tmp(2,49) := "11111111";
			tmp(2,50) := "11111111";
			tmp(2,51) := "11111111";
			tmp(2,52) := "11111111";
			tmp(2,53) := "11111111";
			tmp(2,54) := "11111111";
			tmp(2,55) := "11111111";
			tmp(2,56) := "11111111";
			tmp(2,57) := "11111111";
			tmp(2,58) := "11111111";
			tmp(2,59) := "11111111";
			tmp(2,60) := "11111111";
			tmp(2,61) := "11111111";
			tmp(2,62) := "11111111";
			tmp(2,63) := "11111111";
			tmp(2,64) := "11111111";
			tmp(2,65) := "11111111";
			tmp(2,66) := "11111111";
			tmp(2,67) := "11111111";
			tmp(2,68) := "11111111";
			tmp(2,69) := "11111111";
			tmp(2,70) := "11111111";
			tmp(2,71) := "11111111";
			tmp(2,72) := "11111111";
			tmp(2,73) := "11111111";
			tmp(2,74) := "11111111";
			tmp(2,75) := "11111111";
			tmp(2,76) := "11111111";
			tmp(2,77) := "11111111";
			tmp(2,78) := "11111111";
			tmp(2,79) := "11111111";
			tmp(2,80) := "11111111";
			tmp(3,1) := "11111111";
			tmp(3,2) := "11111111";
			tmp(3,3) := "11111111";
			tmp(3,4) := "11111111";
			tmp(3,5) := "11111111";
			tmp(3,6) := "11111111";
			tmp(3,7) := "11111111";
			tmp(3,8) := "11111111";
			tmp(3,9) := "11111111";
			tmp(3,10) := "11111111";
			tmp(3,11) := "11111111";
			tmp(3,12) := "11111111";
			tmp(3,13) := "11111111";
			tmp(3,14) := "11111111";
			tmp(3,15) := "11111111";
			tmp(3,16) := "11111111";
			tmp(3,17) := "11111111";
			tmp(3,18) := "11111111";
			tmp(3,19) := "11111111";
			tmp(3,20) := "11111111";
			tmp(3,21) := "11111111";
			tmp(3,22) := "11111111";
			tmp(3,23) := "11111111";
			tmp(3,24) := "11111111";
			tmp(3,25) := "11111111";
			tmp(3,26) := "11111111";
			tmp(3,27) := "11111111";
			tmp(3,28) := "11111111";
			tmp(3,29) := "11111111";
			tmp(3,30) := "11111111";
			tmp(3,31) := "11111111";
			tmp(3,32) := "11111111";
			tmp(3,33) := "11111111";
			tmp(3,34) := "11111111";
			tmp(3,35) := "11111111";
			tmp(3,36) := "11111111";
			tmp(3,37) := "11111111";
			tmp(3,38) := "11111111";
			tmp(3,39) := "11111111";
			tmp(3,40) := "11111111";
			tmp(3,41) := "11111111";
			tmp(3,42) := "11111111";
			tmp(3,43) := "11111111";
			tmp(3,44) := "11111111";
			tmp(3,45) := "11111111";
			tmp(3,46) := "11111111";
			tmp(3,47) := "11111111";
			tmp(3,48) := "11111111";
			tmp(3,49) := "11111111";
			tmp(3,50) := "11111111";
			tmp(3,51) := "11111111";
			tmp(3,52) := "11111111";
			tmp(3,53) := "11111111";
			tmp(3,54) := "11111111";
			tmp(3,55) := "11111111";
			tmp(3,56) := "11111111";
			tmp(3,57) := "11111111";
			tmp(3,58) := "11111111";
			tmp(3,59) := "11111111";
			tmp(3,60) := "11111111";
			tmp(3,61) := "11111111";
			tmp(3,62) := "11111111";
			tmp(3,63) := "11111111";
			tmp(3,64) := "11111111";
			tmp(3,65) := "11111111";
			tmp(3,66) := "11111111";
			tmp(3,67) := "11111111";
			tmp(3,68) := "11111111";
			tmp(3,69) := "11111111";
			tmp(3,70) := "11111111";
			tmp(3,71) := "11111111";
			tmp(3,72) := "11111111";
			tmp(3,73) := "11111111";
			tmp(3,74) := "11111111";
			tmp(3,75) := "11111111";
			tmp(3,76) := "11111111";
			tmp(3,77) := "11111111";
			tmp(3,78) := "11111111";
			tmp(3,79) := "11111111";
			tmp(3,80) := "11111111";
			tmp(4,1) := "11111111";
			tmp(4,2) := "11111111";
			tmp(4,3) := "11111111";
			tmp(4,4) := "11111111";
			tmp(4,5) := "11111111";
			tmp(4,6) := "11111111";
			tmp(4,7) := "11111111";
			tmp(4,8) := "11111111";
			tmp(4,9) := "11111111";
			tmp(4,10) := "11111111";
			tmp(4,11) := "11111111";
			tmp(4,12) := "11111111";
			tmp(4,13) := "11111111";
			tmp(4,14) := "11111111";
			tmp(4,15) := "11111111";
			tmp(4,16) := "11111111";
			tmp(4,17) := "11111111";
			tmp(4,18) := "11111111";
			tmp(4,19) := "11111111";
			tmp(4,20) := "11111111";
			tmp(4,21) := "11111111";
			tmp(4,22) := "11111111";
			tmp(4,23) := "11111111";
			tmp(4,24) := "11111111";
			tmp(4,25) := "11111111";
			tmp(4,26) := "11111111";
			tmp(4,27) := "11111111";
			tmp(4,28) := "11111111";
			tmp(4,29) := "11111111";
			tmp(4,30) := "11111111";
			tmp(4,31) := "11111111";
			tmp(4,32) := "11111111";
			tmp(4,33) := "11111111";
			tmp(4,34) := "11111111";
			tmp(4,35) := "11111111";
			tmp(4,36) := "11111111";
			tmp(4,37) := "11111111";
			tmp(4,38) := "11111111";
			tmp(4,39) := "11111111";
			tmp(4,40) := "11111111";
			tmp(4,41) := "11111111";
			tmp(4,42) := "11111111";
			tmp(4,43) := "11111111";
			tmp(4,44) := "11111111";
			tmp(4,45) := "11111111";
			tmp(4,46) := "11111111";
			tmp(4,47) := "11111111";
			tmp(4,48) := "11111111";
			tmp(4,49) := "11111111";
			tmp(4,50) := "11111111";
			tmp(4,51) := "11111111";
			tmp(4,52) := "11111111";
			tmp(4,53) := "11111111";
			tmp(4,54) := "11111111";
			tmp(4,55) := "11111111";
			tmp(4,56) := "11111111";
			tmp(4,57) := "11111111";
			tmp(4,58) := "11111111";
			tmp(4,59) := "11111111";
			tmp(4,60) := "11111111";
			tmp(4,61) := "11111111";
			tmp(4,62) := "11111111";
			tmp(4,63) := "11111111";
			tmp(4,64) := "11111111";
			tmp(4,65) := "11111111";
			tmp(4,66) := "11111111";
			tmp(4,67) := "11111111";
			tmp(4,68) := "11111111";
			tmp(4,69) := "11111111";
			tmp(4,70) := "11111111";
			tmp(4,71) := "11111111";
			tmp(4,72) := "11111111";
			tmp(4,73) := "11111111";
			tmp(4,74) := "11111111";
			tmp(4,75) := "11111111";
			tmp(4,76) := "11111111";
			tmp(4,77) := "11111111";
			tmp(4,78) := "11111111";
			tmp(4,79) := "11111111";
			tmp(4,80) := "11111111";
			tmp(5,1) := "11111111";
			tmp(5,2) := "11111111";
			tmp(5,3) := "11111111";
			tmp(5,4) := "11111111";
			tmp(5,5) := "11111111";
			tmp(5,6) := "11111111";
			tmp(5,7) := "11111111";
			tmp(5,8) := "11111111";
			tmp(5,9) := "11111111";
			tmp(5,10) := "11111111";
			tmp(5,11) := "11111111";
			tmp(5,12) := "11111111";
			tmp(5,13) := "11111111";
			tmp(5,14) := "11111111";
			tmp(5,15) := "11111111";
			tmp(5,16) := "11111111";
			tmp(5,17) := "11111111";
			tmp(5,18) := "11111111";
			tmp(5,19) := "11111111";
			tmp(5,20) := "11111111";
			tmp(5,21) := "11111111";
			tmp(5,22) := "11111111";
			tmp(5,23) := "11111111";
			tmp(5,24) := "11111111";
			tmp(5,25) := "11111111";
			tmp(5,26) := "11111111";
			tmp(5,27) := "11111111";
			tmp(5,28) := "11111111";
			tmp(5,29) := "11111111";
			tmp(5,30) := "11111111";
			tmp(5,31) := "11111111";
			tmp(5,32) := "11111111";
			tmp(5,33) := "11111111";
			tmp(5,34) := "11111111";
			tmp(5,35) := "11111111";
			tmp(5,36) := "11111111";
			tmp(5,37) := "11111111";
			tmp(5,38) := "11111111";
			tmp(5,39) := "11111111";
			tmp(5,40) := "11111111";
			tmp(5,41) := "11111111";
			tmp(5,42) := "11111111";
			tmp(5,43) := "11111111";
			tmp(5,44) := "11111111";
			tmp(5,45) := "11111111";
			tmp(5,46) := "11111111";
			tmp(5,47) := "11111111";
			tmp(5,48) := "11111111";
			tmp(5,49) := "11111111";
			tmp(5,50) := "11111111";
			tmp(5,51) := "11111111";
			tmp(5,52) := "11111111";
			tmp(5,53) := "11111111";
			tmp(5,54) := "11111111";
			tmp(5,55) := "11111111";
			tmp(5,56) := "11111111";
			tmp(5,57) := "11111111";
			tmp(5,58) := "11111111";
			tmp(5,59) := "11111111";
			tmp(5,60) := "11111111";
			tmp(5,61) := "11111111";
			tmp(5,62) := "11111111";
			tmp(5,63) := "11111111";
			tmp(5,64) := "11111111";
			tmp(5,65) := "11111111";
			tmp(5,66) := "11111111";
			tmp(5,67) := "11111111";
			tmp(5,68) := "11111111";
			tmp(5,69) := "11111111";
			tmp(5,70) := "11111111";
			tmp(5,71) := "11111111";
			tmp(5,72) := "11111111";
			tmp(5,73) := "11111111";
			tmp(5,74) := "11111111";
			tmp(5,75) := "11111111";
			tmp(5,76) := "11111111";
			tmp(5,77) := "11111111";
			tmp(5,78) := "11111111";
			tmp(5,79) := "11111111";
			tmp(5,80) := "11111111";
			tmp(6,1) := "11111111";
			tmp(6,2) := "11111111";
			tmp(6,3) := "11111111";
			tmp(6,4) := "11111111";
			tmp(6,5) := "11111111";
			tmp(6,6) := "11111111";
			tmp(6,7) := "11111111";
			tmp(6,8) := "11111111";
			tmp(6,9) := "11111111";
			tmp(6,10) := "11111111";
			tmp(6,11) := "11111111";
			tmp(6,12) := "11111111";
			tmp(6,13) := "11111111";
			tmp(6,14) := "11111111";
			tmp(6,15) := "11111111";
			tmp(6,16) := "11111111";
			tmp(6,17) := "11111111";
			tmp(6,18) := "11111111";
			tmp(6,19) := "11111111";
			tmp(6,20) := "11111111";
			tmp(6,21) := "11111111";
			tmp(6,22) := "11111111";
			tmp(6,23) := "11111111";
			tmp(6,24) := "11111111";
			tmp(6,25) := "11111111";
			tmp(6,26) := "11111111";
			tmp(6,27) := "11111111";
			tmp(6,28) := "11111111";
			tmp(6,29) := "11111111";
			tmp(6,30) := "11111111";
			tmp(6,31) := "11111111";
			tmp(6,32) := "11111111";
			tmp(6,33) := "11111111";
			tmp(6,34) := "11111111";
			tmp(6,35) := "11111111";
			tmp(6,36) := "11111111";
			tmp(6,37) := "11111111";
			tmp(6,38) := "11111111";
			tmp(6,39) := "11111111";
			tmp(6,40) := "11111111";
			tmp(6,41) := "11111111";
			tmp(6,42) := "11111111";
			tmp(6,43) := "11111111";
			tmp(6,44) := "11111111";
			tmp(6,45) := "11111111";
			tmp(6,46) := "11111111";
			tmp(6,47) := "11111111";
			tmp(6,48) := "11111111";
			tmp(6,49) := "11111111";
			tmp(6,50) := "11111111";
			tmp(6,51) := "11111111";
			tmp(6,52) := "11111111";
			tmp(6,53) := "11111111";
			tmp(6,54) := "11111111";
			tmp(6,55) := "11111111";
			tmp(6,56) := "11111111";
			tmp(6,57) := "11111111";
			tmp(6,58) := "11111111";
			tmp(6,59) := "11111111";
			tmp(6,60) := "11111111";
			tmp(6,61) := "11111111";
			tmp(6,62) := "11111111";
			tmp(6,63) := "11111111";
			tmp(6,64) := "11111111";
			tmp(6,65) := "11111111";
			tmp(6,66) := "11111111";
			tmp(6,67) := "11111111";
			tmp(6,68) := "11111111";
			tmp(6,69) := "11111111";
			tmp(6,70) := "11111111";
			tmp(6,71) := "11111111";
			tmp(6,72) := "11111111";
			tmp(6,73) := "11111111";
			tmp(6,74) := "11111111";
			tmp(6,75) := "11111111";
			tmp(6,76) := "11111111";
			tmp(6,77) := "11111111";
			tmp(6,78) := "11111111";
			tmp(6,79) := "11111111";
			tmp(6,80) := "11111111";
			tmp(7,1) := "11111111";
			tmp(7,2) := "11111111";
			tmp(7,3) := "11111111";
			tmp(7,4) := "11111111";
			tmp(7,5) := "11111111";
			tmp(7,6) := "11111111";
			tmp(7,7) := "11111111";
			tmp(7,8) := "11111111";
			tmp(7,9) := "11111111";
			tmp(7,10) := "11111111";
			tmp(7,11) := "11111111";
			tmp(7,12) := "11111111";
			tmp(7,13) := "11111111";
			tmp(7,14) := "11111111";
			tmp(7,15) := "11111111";
			tmp(7,16) := "11111111";
			tmp(7,17) := "11111111";
			tmp(7,18) := "11111111";
			tmp(7,19) := "11111111";
			tmp(7,20) := "11111111";
			tmp(7,21) := "11111111";
			tmp(7,22) := "11111111";
			tmp(7,23) := "11111111";
			tmp(7,24) := "11111111";
			tmp(7,25) := "11111111";
			tmp(7,26) := "11111111";
			tmp(7,27) := "11111111";
			tmp(7,28) := "11111111";
			tmp(7,29) := "11111111";
			tmp(7,30) := "11111111";
			tmp(7,31) := "11111111";
			tmp(7,32) := "11111111";
			tmp(7,33) := "11111111";
			tmp(7,34) := "11111111";
			tmp(7,35) := "11111111";
			tmp(7,36) := "11111111";
			tmp(7,37) := "11111111";
			tmp(7,38) := "11111111";
			tmp(7,39) := "11111111";
			tmp(7,40) := "11111111";
			tmp(7,41) := "11111111";
			tmp(7,42) := "11111111";
			tmp(7,43) := "11111111";
			tmp(7,44) := "11111111";
			tmp(7,45) := "11111111";
			tmp(7,46) := "11111111";
			tmp(7,47) := "11111111";
			tmp(7,48) := "11111111";
			tmp(7,49) := "11111111";
			tmp(7,50) := "11111111";
			tmp(7,51) := "11111111";
			tmp(7,52) := "11111111";
			tmp(7,53) := "11111111";
			tmp(7,54) := "11111111";
			tmp(7,55) := "11111111";
			tmp(7,56) := "11111111";
			tmp(7,57) := "11111111";
			tmp(7,58) := "11111111";
			tmp(7,59) := "11111111";
			tmp(7,60) := "11111111";
			tmp(7,61) := "11111111";
			tmp(7,62) := "11111111";
			tmp(7,63) := "11111111";
			tmp(7,64) := "11111111";
			tmp(7,65) := "11111111";
			tmp(7,66) := "11111111";
			tmp(7,67) := "11111111";
			tmp(7,68) := "11111111";
			tmp(7,69) := "11111111";
			tmp(7,70) := "11111111";
			tmp(7,71) := "11111111";
			tmp(7,72) := "11111111";
			tmp(7,73) := "11111111";
			tmp(7,74) := "11111111";
			tmp(7,75) := "11111111";
			tmp(7,76) := "11111111";
			tmp(7,77) := "11111111";
			tmp(7,78) := "11111111";
			tmp(7,79) := "11111111";
			tmp(7,80) := "11111111";
			tmp(8,1) := "11111111";
			tmp(8,2) := "11111111";
			tmp(8,3) := "11111111";
			tmp(8,4) := "11111111";
			tmp(8,5) := "11111111";
			tmp(8,6) := "11111111";
			tmp(8,7) := "11111111";
			tmp(8,8) := "11111111";
			tmp(8,9) := "11111111";
			tmp(8,10) := "11111111";
			tmp(8,11) := "11111111";
			tmp(8,12) := "11111111";
			tmp(8,13) := "11111111";
			tmp(8,14) := "11111111";
			tmp(8,15) := "11111111";
			tmp(8,16) := "11111111";
			tmp(8,17) := "11111111";
			tmp(8,18) := "11111111";
			tmp(8,19) := "11111111";
			tmp(8,20) := "11111111";
			tmp(8,21) := "11111111";
			tmp(8,22) := "11111111";
			tmp(8,23) := "11111111";
			tmp(8,24) := "11111111";
			tmp(8,25) := "11111111";
			tmp(8,26) := "11111111";
			tmp(8,27) := "11111111";
			tmp(8,28) := "11111111";
			tmp(8,29) := "11111111";
			tmp(8,30) := "11111111";
			tmp(8,31) := "11111111";
			tmp(8,32) := "11111111";
			tmp(8,33) := "11111111";
			tmp(8,34) := "11111111";
			tmp(8,35) := "11111111";
			tmp(8,36) := "11111111";
			tmp(8,37) := "11111111";
			tmp(8,38) := "11111111";
			tmp(8,39) := "11111111";
			tmp(8,40) := "11111111";
			tmp(8,41) := "11111111";
			tmp(8,42) := "11111111";
			tmp(8,43) := "11111111";
			tmp(8,44) := "11111111";
			tmp(8,45) := "11111111";
			tmp(8,46) := "11111111";
			tmp(8,47) := "11111111";
			tmp(8,48) := "11111111";
			tmp(8,49) := "11111111";
			tmp(8,50) := "11111111";
			tmp(8,51) := "11111111";
			tmp(8,52) := "11111111";
			tmp(8,53) := "11111111";
			tmp(8,54) := "11111111";
			tmp(8,55) := "11111111";
			tmp(8,56) := "11111111";
			tmp(8,57) := "11111111";
			tmp(8,58) := "11111111";
			tmp(8,59) := "11111111";
			tmp(8,60) := "11111111";
			tmp(8,61) := "11111111";
			tmp(8,62) := "11111111";
			tmp(8,63) := "11111111";
			tmp(8,64) := "11111111";
			tmp(8,65) := "11111111";
			tmp(8,66) := "11111111";
			tmp(8,67) := "11111111";
			tmp(8,68) := "11111111";
			tmp(8,69) := "11111111";
			tmp(8,70) := "11111111";
			tmp(8,71) := "11111111";
			tmp(8,72) := "11111111";
			tmp(8,73) := "11111111";
			tmp(8,74) := "11111111";
			tmp(8,75) := "11111111";
			tmp(8,76) := "11111111";
			tmp(8,77) := "11111111";
			tmp(8,78) := "11111111";
			tmp(8,79) := "11111111";
			tmp(8,80) := "11111111";
			tmp(9,1) := "11111111";
			tmp(9,2) := "11111111";
			tmp(9,3) := "11111111";
			tmp(9,4) := "11111111";
			tmp(9,5) := "11111111";
			tmp(9,6) := "11111111";
			tmp(9,7) := "11111111";
			tmp(9,8) := "11111111";
			tmp(9,9) := "11111111";
			tmp(9,10) := "11111111";
			tmp(9,11) := "11111111";
			tmp(9,12) := "11111111";
			tmp(9,13) := "11111111";
			tmp(9,14) := "11111111";
			tmp(9,15) := "11111111";
			tmp(9,16) := "11111111";
			tmp(9,17) := "11111111";
			tmp(9,18) := "11111111";
			tmp(9,19) := "11111111";
			tmp(9,20) := "11111111";
			tmp(9,21) := "11111111";
			tmp(9,22) := "11111111";
			tmp(9,23) := "11111111";
			tmp(9,24) := "11111111";
			tmp(9,25) := "11111111";
			tmp(9,26) := "11111111";
			tmp(9,27) := "11111111";
			tmp(9,28) := "11111111";
			tmp(9,29) := "11111111";
			tmp(9,30) := "11111111";
			tmp(9,31) := "11111111";
			tmp(9,32) := "11111111";
			tmp(9,33) := "11111111";
			tmp(9,34) := "11111011";
			tmp(9,35) := "11111111";
			tmp(9,36) := "11111111";
			tmp(9,37) := "11111111";
			tmp(9,38) := "11111110";
			tmp(9,39) := "11111110";
			tmp(9,40) := "11111111";
			tmp(9,41) := "11111111";
			tmp(9,42) := "11111110";
			tmp(9,43) := "11111111";
			tmp(9,44) := "11111110";
			tmp(9,45) := "11111111";
			tmp(9,46) := "11111011";
			tmp(9,47) := "11111110";
			tmp(9,48) := "11111111";
			tmp(9,49) := "11111110";
			tmp(9,50) := "11111111";
			tmp(9,51) := "11111100";
			tmp(9,52) := "11111001";
			tmp(9,53) := "11111101";
			tmp(9,54) := "11110010";
			tmp(9,55) := "11110001";
			tmp(9,56) := "11111100";
			tmp(9,57) := "11111011";
			tmp(9,58) := "11111011";
			tmp(9,59) := "11111100";
			tmp(9,60) := "11111111";
			tmp(9,61) := "11111111";
			tmp(9,62) := "11111111";
			tmp(9,63) := "11111110";
			tmp(9,64) := "11111111";
			tmp(9,65) := "11111111";
			tmp(9,66) := "11111110";
			tmp(9,67) := "11111110";
			tmp(9,68) := "11111111";
			tmp(9,69) := "11111111";
			tmp(9,70) := "11111111";
			tmp(9,71) := "11111110";
			tmp(9,72) := "11111110";
			tmp(9,73) := "11111100";
			tmp(9,74) := "11111100";
			tmp(9,75) := "11111111";
			tmp(9,76) := "11111110";
			tmp(9,77) := "11111010";
			tmp(9,78) := "11111100";
			tmp(9,79) := "11111111";
			tmp(9,80) := "11111111";
			tmp(10,1) := "11111111";
			tmp(10,2) := "11111111";
			tmp(10,3) := "11111111";
			tmp(10,4) := "11111111";
			tmp(10,5) := "11111111";
			tmp(10,6) := "11111111";
			tmp(10,7) := "11111111";
			tmp(10,8) := "11111111";
			tmp(10,9) := "11111111";
			tmp(10,10) := "11111111";
			tmp(10,11) := "11111111";
			tmp(10,12) := "11111111";
			tmp(10,13) := "11111111";
			tmp(10,14) := "11111111";
			tmp(10,15) := "11111111";
			tmp(10,16) := "11111111";
			tmp(10,17) := "11111111";
			tmp(10,18) := "11111111";
			tmp(10,19) := "11111111";
			tmp(10,20) := "11111111";
			tmp(10,21) := "11111111";
			tmp(10,22) := "11111111";
			tmp(10,23) := "11111111";
			tmp(10,24) := "11111111";
			tmp(10,25) := "11111111";
			tmp(10,26) := "11111111";
			tmp(10,27) := "11111111";
			tmp(10,28) := "11111111";
			tmp(10,29) := "11111111";
			tmp(10,30) := "11111111";
			tmp(10,31) := "11111111";
			tmp(10,32) := "11111111";
			tmp(10,33) := "11111110";
			tmp(10,34) := "11111111";
			tmp(10,35) := "11111101";
			tmp(10,36) := "11111001";
			tmp(10,37) := "11111100";
			tmp(10,38) := "11111100";
			tmp(10,39) := "11111010";
			tmp(10,40) := "11111111";
			tmp(10,41) := "11111011";
			tmp(10,42) := "11111110";
			tmp(10,43) := "11111100";
			tmp(10,44) := "11111111";
			tmp(10,45) := "11111111";
			tmp(10,46) := "11111011";
			tmp(10,47) := "11111111";
			tmp(10,48) := "11111101";
			tmp(10,49) := "11111101";
			tmp(10,50) := "11110110";
			tmp(10,51) := "11101000";
			tmp(10,52) := "11110001";
			tmp(10,53) := "11010110";
			tmp(10,54) := "11000100";
			tmp(10,55) := "11001001";
			tmp(10,56) := "11001110";
			tmp(10,57) := "11010010";
			tmp(10,58) := "10111110";
			tmp(10,59) := "11000011";
			tmp(10,60) := "11001011";
			tmp(10,61) := "11011101";
			tmp(10,62) := "11110101";
			tmp(10,63) := "11111001";
			tmp(10,64) := "11111011";
			tmp(10,65) := "11111011";
			tmp(10,66) := "11111111";
			tmp(10,67) := "11111101";
			tmp(10,68) := "11111100";
			tmp(10,69) := "11111110";
			tmp(10,70) := "11111111";
			tmp(10,71) := "11111111";
			tmp(10,72) := "11111111";
			tmp(10,73) := "11111111";
			tmp(10,74) := "11111111";
			tmp(10,75) := "11111110";
			tmp(10,76) := "11111111";
			tmp(10,77) := "11111110";
			tmp(10,78) := "11111101";
			tmp(10,79) := "11111101";
			tmp(10,80) := "11111111";
			tmp(11,1) := "11111111";
			tmp(11,2) := "11111111";
			tmp(11,3) := "11111111";
			tmp(11,4) := "11111111";
			tmp(11,5) := "11111111";
			tmp(11,6) := "11111111";
			tmp(11,7) := "11111111";
			tmp(11,8) := "11111111";
			tmp(11,9) := "11111111";
			tmp(11,10) := "11111111";
			tmp(11,11) := "11111111";
			tmp(11,12) := "11111111";
			tmp(11,13) := "11111111";
			tmp(11,14) := "11111111";
			tmp(11,15) := "11111111";
			tmp(11,16) := "11111111";
			tmp(11,17) := "11111111";
			tmp(11,18) := "11111111";
			tmp(11,19) := "11111111";
			tmp(11,20) := "11111111";
			tmp(11,21) := "11111111";
			tmp(11,22) := "11111111";
			tmp(11,23) := "11111111";
			tmp(11,24) := "11111111";
			tmp(11,25) := "11111111";
			tmp(11,26) := "11111111";
			tmp(11,27) := "11111111";
			tmp(11,28) := "11111111";
			tmp(11,29) := "11111111";
			tmp(11,30) := "11111111";
			tmp(11,31) := "11111111";
			tmp(11,32) := "11111111";
			tmp(11,33) := "11111111";
			tmp(11,34) := "11110111";
			tmp(11,35) := "11111011";
			tmp(11,36) := "11111111";
			tmp(11,37) := "11111111";
			tmp(11,38) := "11111111";
			tmp(11,39) := "11111111";
			tmp(11,40) := "11111101";
			tmp(11,41) := "11111111";
			tmp(11,42) := "11111111";
			tmp(11,43) := "11111111";
			tmp(11,44) := "11111111";
			tmp(11,45) := "11111010";
			tmp(11,46) := "11111100";
			tmp(11,47) := "11110000";
			tmp(11,48) := "11110010";
			tmp(11,49) := "11101001";
			tmp(11,50) := "11011000";
			tmp(11,51) := "11011111";
			tmp(11,52) := "11101000";
			tmp(11,53) := "11010111";
			tmp(11,54) := "10111011";
			tmp(11,55) := "11000011";
			tmp(11,56) := "11001010";
			tmp(11,57) := "11000100";
			tmp(11,58) := "10111010";
			tmp(11,59) := "10110000";
			tmp(11,60) := "10111010";
			tmp(11,61) := "10110110";
			tmp(11,62) := "10101101";
			tmp(11,63) := "11000000";
			tmp(11,64) := "11001010";
			tmp(11,65) := "11011001";
			tmp(11,66) := "11101111";
			tmp(11,67) := "11111111";
			tmp(11,68) := "11111110";
			tmp(11,69) := "11111100";
			tmp(11,70) := "11111100";
			tmp(11,71) := "11111111";
			tmp(11,72) := "11111110";
			tmp(11,73) := "11111110";
			tmp(11,74) := "11111111";
			tmp(11,75) := "11111111";
			tmp(11,76) := "11111111";
			tmp(11,77) := "11111110";
			tmp(11,78) := "11111110";
			tmp(11,79) := "11111111";
			tmp(11,80) := "11111110";
			tmp(12,1) := "11111111";
			tmp(12,2) := "11111111";
			tmp(12,3) := "11111111";
			tmp(12,4) := "11111111";
			tmp(12,5) := "11111111";
			tmp(12,6) := "11111111";
			tmp(12,7) := "11111111";
			tmp(12,8) := "11111111";
			tmp(12,9) := "11111111";
			tmp(12,10) := "11111111";
			tmp(12,11) := "11111111";
			tmp(12,12) := "11111111";
			tmp(12,13) := "11111111";
			tmp(12,14) := "11111111";
			tmp(12,15) := "11111111";
			tmp(12,16) := "11111111";
			tmp(12,17) := "11111111";
			tmp(12,18) := "11111111";
			tmp(12,19) := "11111111";
			tmp(12,20) := "11111111";
			tmp(12,21) := "11111111";
			tmp(12,22) := "11111111";
			tmp(12,23) := "11111111";
			tmp(12,24) := "11111111";
			tmp(12,25) := "11111111";
			tmp(12,26) := "11111111";
			tmp(12,27) := "11111111";
			tmp(12,28) := "11111111";
			tmp(12,29) := "11111111";
			tmp(12,30) := "11111111";
			tmp(12,31) := "11111111";
			tmp(12,32) := "11111111";
			tmp(12,33) := "11111111";
			tmp(12,34) := "11111111";
			tmp(12,35) := "11111110";
			tmp(12,36) := "11111100";
			tmp(12,37) := "11111111";
			tmp(12,38) := "11111101";
			tmp(12,39) := "11111110";
			tmp(12,40) := "11111110";
			tmp(12,41) := "11111110";
			tmp(12,42) := "11111110";
			tmp(12,43) := "11111111";
			tmp(12,44) := "11101110";
			tmp(12,45) := "11101011";
			tmp(12,46) := "11011010";
			tmp(12,47) := "11010101";
			tmp(12,48) := "11011100";
			tmp(12,49) := "11010111";
			tmp(12,50) := "11010000";
			tmp(12,51) := "11011100";
			tmp(12,52) := "11001111";
			tmp(12,53) := "11000111";
			tmp(12,54) := "10111000";
			tmp(12,55) := "10101110";
			tmp(12,56) := "10111011";
			tmp(12,57) := "10110111";
			tmp(12,58) := "10101111";
			tmp(12,59) := "10101100";
			tmp(12,60) := "10110110";
			tmp(12,61) := "10101111";
			tmp(12,62) := "10011100";
			tmp(12,63) := "10100011";
			tmp(12,64) := "10101000";
			tmp(12,65) := "10100000";
			tmp(12,66) := "10100101";
			tmp(12,67) := "11000110";
			tmp(12,68) := "11101001";
			tmp(12,69) := "11111111";
			tmp(12,70) := "11111100";
			tmp(12,71) := "11111110";
			tmp(12,72) := "11111111";
			tmp(12,73) := "11111111";
			tmp(12,74) := "11111101";
			tmp(12,75) := "11111111";
			tmp(12,76) := "11111111";
			tmp(12,77) := "11111111";
			tmp(12,78) := "11111111";
			tmp(12,79) := "11111111";
			tmp(12,80) := "11111111";
			tmp(13,1) := "11111111";
			tmp(13,2) := "11111111";
			tmp(13,3) := "11111111";
			tmp(13,4) := "11111111";
			tmp(13,5) := "11111111";
			tmp(13,6) := "11111111";
			tmp(13,7) := "11111111";
			tmp(13,8) := "11111111";
			tmp(13,9) := "11111111";
			tmp(13,10) := "11111111";
			tmp(13,11) := "11111111";
			tmp(13,12) := "11111111";
			tmp(13,13) := "11111111";
			tmp(13,14) := "11111111";
			tmp(13,15) := "11111111";
			tmp(13,16) := "11111111";
			tmp(13,17) := "11111111";
			tmp(13,18) := "11111111";
			tmp(13,19) := "11111111";
			tmp(13,20) := "11111111";
			tmp(13,21) := "11111111";
			tmp(13,22) := "11111111";
			tmp(13,23) := "11111111";
			tmp(13,24) := "11111111";
			tmp(13,25) := "11111111";
			tmp(13,26) := "11111111";
			tmp(13,27) := "11111111";
			tmp(13,28) := "11111111";
			tmp(13,29) := "11111111";
			tmp(13,30) := "11111111";
			tmp(13,31) := "11111111";
			tmp(13,32) := "11111111";
			tmp(13,33) := "11111110";
			tmp(13,34) := "11111100";
			tmp(13,35) := "11111011";
			tmp(13,36) := "11111111";
			tmp(13,37) := "11111111";
			tmp(13,38) := "11111000";
			tmp(13,39) := "11111101";
			tmp(13,40) := "11111001";
			tmp(13,41) := "11110110";
			tmp(13,42) := "11110010";
			tmp(13,43) := "11100010";
			tmp(13,44) := "11010111";
			tmp(13,45) := "11011110";
			tmp(13,46) := "11001110";
			tmp(13,47) := "11010101";
			tmp(13,48) := "11011000";
			tmp(13,49) := "11010001";
			tmp(13,50) := "11000110";
			tmp(13,51) := "11000100";
			tmp(13,52) := "11000111";
			tmp(13,53) := "10111010";
			tmp(13,54) := "10100001";
			tmp(13,55) := "10100110";
			tmp(13,56) := "10110110";
			tmp(13,57) := "10110111";
			tmp(13,58) := "10010111";
			tmp(13,59) := "10011011";
			tmp(13,60) := "10101011";
			tmp(13,61) := "10100111";
			tmp(13,62) := "10011011";
			tmp(13,63) := "10011000";
			tmp(13,64) := "10100001";
			tmp(13,65) := "10011110";
			tmp(13,66) := "10011011";
			tmp(13,67) := "10100111";
			tmp(13,68) := "10011001";
			tmp(13,69) := "11011011";
			tmp(13,70) := "11111111";
			tmp(13,71) := "11111101";
			tmp(13,72) := "11111110";
			tmp(13,73) := "11111110";
			tmp(13,74) := "11111110";
			tmp(13,75) := "11111110";
			tmp(13,76) := "11111101";
			tmp(13,77) := "11111111";
			tmp(13,78) := "11111111";
			tmp(13,79) := "11111100";
			tmp(13,80) := "11111111";
			tmp(14,1) := "11111111";
			tmp(14,2) := "11111111";
			tmp(14,3) := "11111111";
			tmp(14,4) := "11111111";
			tmp(14,5) := "11111111";
			tmp(14,6) := "11111111";
			tmp(14,7) := "11111111";
			tmp(14,8) := "11111111";
			tmp(14,9) := "11111111";
			tmp(14,10) := "11111111";
			tmp(14,11) := "11111111";
			tmp(14,12) := "11111111";
			tmp(14,13) := "11111111";
			tmp(14,14) := "11111111";
			tmp(14,15) := "11111111";
			tmp(14,16) := "11111111";
			tmp(14,17) := "11111111";
			tmp(14,18) := "11111111";
			tmp(14,19) := "11111111";
			tmp(14,20) := "11111111";
			tmp(14,21) := "11111111";
			tmp(14,22) := "11111111";
			tmp(14,23) := "11111111";
			tmp(14,24) := "11111111";
			tmp(14,25) := "11111111";
			tmp(14,26) := "11111111";
			tmp(14,27) := "11111111";
			tmp(14,28) := "11111111";
			tmp(14,29) := "11111111";
			tmp(14,30) := "11111111";
			tmp(14,31) := "11111111";
			tmp(14,32) := "11111111";
			tmp(14,33) := "11111110";
			tmp(14,34) := "11111110";
			tmp(14,35) := "11111111";
			tmp(14,36) := "11111111";
			tmp(14,37) := "11111000";
			tmp(14,38) := "11111111";
			tmp(14,39) := "11101010";
			tmp(14,40) := "11100101";
			tmp(14,41) := "11100100";
			tmp(14,42) := "11100001";
			tmp(14,43) := "11100000";
			tmp(14,44) := "11010010";
			tmp(14,45) := "11001000";
			tmp(14,46) := "10111111";
			tmp(14,47) := "10110110";
			tmp(14,48) := "11000100";
			tmp(14,49) := "11000011";
			tmp(14,50) := "10111101";
			tmp(14,51) := "10111010";
			tmp(14,52) := "10111011";
			tmp(14,53) := "10101100";
			tmp(14,54) := "10100001";
			tmp(14,55) := "10100100";
			tmp(14,56) := "10101110";
			tmp(14,57) := "10100011";
			tmp(14,58) := "10010101";
			tmp(14,59) := "10011010";
			tmp(14,60) := "10100011";
			tmp(14,61) := "10011110";
			tmp(14,62) := "10010100";
			tmp(14,63) := "10010110";
			tmp(14,64) := "10010001";
			tmp(14,65) := "10001111";
			tmp(14,66) := "10010100";
			tmp(14,67) := "10010110";
			tmp(14,68) := "10010110";
			tmp(14,69) := "10011100";
			tmp(14,70) := "11001001";
			tmp(14,71) := "11101111";
			tmp(14,72) := "11111110";
			tmp(14,73) := "11111111";
			tmp(14,74) := "11111100";
			tmp(14,75) := "11111100";
			tmp(14,76) := "11111101";
			tmp(14,77) := "11111110";
			tmp(14,78) := "11111111";
			tmp(14,79) := "11111111";
			tmp(14,80) := "11111110";
			tmp(15,1) := "11111111";
			tmp(15,2) := "11111111";
			tmp(15,3) := "11111111";
			tmp(15,4) := "11111111";
			tmp(15,5) := "11111111";
			tmp(15,6) := "11111111";
			tmp(15,7) := "11111111";
			tmp(15,8) := "11111111";
			tmp(15,9) := "11111111";
			tmp(15,10) := "11111111";
			tmp(15,11) := "11111111";
			tmp(15,12) := "11111111";
			tmp(15,13) := "11111111";
			tmp(15,14) := "11111111";
			tmp(15,15) := "11111111";
			tmp(15,16) := "11111111";
			tmp(15,17) := "11111111";
			tmp(15,18) := "11111111";
			tmp(15,19) := "11111111";
			tmp(15,20) := "11111111";
			tmp(15,21) := "11111111";
			tmp(15,22) := "11111111";
			tmp(15,23) := "11111111";
			tmp(15,24) := "11111111";
			tmp(15,25) := "11111111";
			tmp(15,26) := "11111111";
			tmp(15,27) := "11111111";
			tmp(15,28) := "11111111";
			tmp(15,29) := "11111111";
			tmp(15,30) := "11111111";
			tmp(15,31) := "11111111";
			tmp(15,32) := "11111111";
			tmp(15,33) := "11111110";
			tmp(15,34) := "11111110";
			tmp(15,35) := "11111010";
			tmp(15,36) := "11111101";
			tmp(15,37) := "11101111";
			tmp(15,38) := "11100011";
			tmp(15,39) := "11011010";
			tmp(15,40) := "11010110";
			tmp(15,41) := "11001101";
			tmp(15,42) := "11010011";
			tmp(15,43) := "11010110";
			tmp(15,44) := "11010010";
			tmp(15,45) := "11001011";
			tmp(15,46) := "10110111";
			tmp(15,47) := "11000010";
			tmp(15,48) := "11000110";
			tmp(15,49) := "11000000";
			tmp(15,50) := "10110100";
			tmp(15,51) := "10111011";
			tmp(15,52) := "10110011";
			tmp(15,53) := "10101010";
			tmp(15,54) := "10100101";
			tmp(15,55) := "10100110";
			tmp(15,56) := "10100111";
			tmp(15,57) := "10011110";
			tmp(15,58) := "10010101";
			tmp(15,59) := "10011101";
			tmp(15,60) := "10100010";
			tmp(15,61) := "10010111";
			tmp(15,62) := "10000111";
			tmp(15,63) := "10000110";
			tmp(15,64) := "10000110";
			tmp(15,65) := "10000010";
			tmp(15,66) := "10000001";
			tmp(15,67) := "10000010";
			tmp(15,68) := "10001000";
			tmp(15,69) := "10010101";
			tmp(15,70) := "10001100";
			tmp(15,71) := "10111011";
			tmp(15,72) := "11101101";
			tmp(15,73) := "11111111";
			tmp(15,74) := "11111111";
			tmp(15,75) := "11111111";
			tmp(15,76) := "11111110";
			tmp(15,77) := "11111111";
			tmp(15,78) := "11111101";
			tmp(15,79) := "11111111";
			tmp(15,80) := "11111111";
			tmp(16,1) := "11111111";
			tmp(16,2) := "11111111";
			tmp(16,3) := "11111111";
			tmp(16,4) := "11111111";
			tmp(16,5) := "11111111";
			tmp(16,6) := "11111111";
			tmp(16,7) := "11111111";
			tmp(16,8) := "11111111";
			tmp(16,9) := "11111111";
			tmp(16,10) := "11111111";
			tmp(16,11) := "11111111";
			tmp(16,12) := "11111111";
			tmp(16,13) := "11111111";
			tmp(16,14) := "11111111";
			tmp(16,15) := "11111111";
			tmp(16,16) := "11111111";
			tmp(16,17) := "11111111";
			tmp(16,18) := "11111111";
			tmp(16,19) := "11111111";
			tmp(16,20) := "11111111";
			tmp(16,21) := "11111111";
			tmp(16,22) := "11111111";
			tmp(16,23) := "11111111";
			tmp(16,24) := "11111111";
			tmp(16,25) := "11111111";
			tmp(16,26) := "11111111";
			tmp(16,27) := "11111111";
			tmp(16,28) := "11111111";
			tmp(16,29) := "11111111";
			tmp(16,30) := "11111111";
			tmp(16,31) := "11111111";
			tmp(16,32) := "11111111";
			tmp(16,33) := "11111010";
			tmp(16,34) := "11110101";
			tmp(16,35) := "11110011";
			tmp(16,36) := "11100011";
			tmp(16,37) := "11110110";
			tmp(16,38) := "11101100";
			tmp(16,39) := "11010001";
			tmp(16,40) := "11001010";
			tmp(16,41) := "11000000";
			tmp(16,42) := "11001010";
			tmp(16,43) := "11001010";
			tmp(16,44) := "11001110";
			tmp(16,45) := "10111100";
			tmp(16,46) := "10101111";
			tmp(16,47) := "10110001";
			tmp(16,48) := "10111001";
			tmp(16,49) := "10101100";
			tmp(16,50) := "10100110";
			tmp(16,51) := "10110010";
			tmp(16,52) := "10110010";
			tmp(16,53) := "10100001";
			tmp(16,54) := "10011110";
			tmp(16,55) := "10010001";
			tmp(16,56) := "10010111";
			tmp(16,57) := "10001110";
			tmp(16,58) := "10000100";
			tmp(16,59) := "10001110";
			tmp(16,60) := "10010011";
			tmp(16,61) := "10000111";
			tmp(16,62) := "10000000";
			tmp(16,63) := "10000101";
			tmp(16,64) := "01111110";
			tmp(16,65) := "01111101";
			tmp(16,66) := "01111111";
			tmp(16,67) := "01110010";
			tmp(16,68) := "01111000";
			tmp(16,69) := "10000001";
			tmp(16,70) := "01111110";
			tmp(16,71) := "10001011";
			tmp(16,72) := "10011010";
			tmp(16,73) := "10101110";
			tmp(16,74) := "11101110";
			tmp(16,75) := "11111111";
			tmp(16,76) := "11111101";
			tmp(16,77) := "11111111";
			tmp(16,78) := "11111110";
			tmp(16,79) := "11111110";
			tmp(16,80) := "11111110";
			tmp(17,1) := "11111111";
			tmp(17,2) := "11111111";
			tmp(17,3) := "11111111";
			tmp(17,4) := "11111111";
			tmp(17,5) := "11111111";
			tmp(17,6) := "11111111";
			tmp(17,7) := "11111111";
			tmp(17,8) := "11111111";
			tmp(17,9) := "11111111";
			tmp(17,10) := "11111111";
			tmp(17,11) := "11111111";
			tmp(17,12) := "11111111";
			tmp(17,13) := "11111111";
			tmp(17,14) := "11111111";
			tmp(17,15) := "11111111";
			tmp(17,16) := "11111111";
			tmp(17,17) := "11111110";
			tmp(17,18) := "11111110";
			tmp(17,19) := "11111111";
			tmp(17,20) := "11111111";
			tmp(17,21) := "11111111";
			tmp(17,22) := "11111110";
			tmp(17,23) := "11111111";
			tmp(17,24) := "11111111";
			tmp(17,25) := "11111111";
			tmp(17,26) := "11111111";
			tmp(17,27) := "11111111";
			tmp(17,28) := "11111000";
			tmp(17,29) := "11111110";
			tmp(17,30) := "11111111";
			tmp(17,31) := "11111101";
			tmp(17,32) := "11111000";
			tmp(17,33) := "11101111";
			tmp(17,34) := "11101010";
			tmp(17,35) := "11100100";
			tmp(17,36) := "11100011";
			tmp(17,37) := "11100000";
			tmp(17,38) := "11011011";
			tmp(17,39) := "11000000";
			tmp(17,40) := "11000100";
			tmp(17,41) := "11000011";
			tmp(17,42) := "11000000";
			tmp(17,43) := "11001000";
			tmp(17,44) := "11001000";
			tmp(17,45) := "10111101";
			tmp(17,46) := "10100011";
			tmp(17,47) := "10101101";
			tmp(17,48) := "10101100";
			tmp(17,49) := "10011111";
			tmp(17,50) := "10011011";
			tmp(17,51) := "10110011";
			tmp(17,52) := "10101010";
			tmp(17,53) := "10011011";
			tmp(17,54) := "10001101";
			tmp(17,55) := "10001010";
			tmp(17,56) := "10001011";
			tmp(17,57) := "10000001";
			tmp(17,58) := "01111110";
			tmp(17,59) := "10000010";
			tmp(17,60) := "10000010";
			tmp(17,61) := "01111100";
			tmp(17,62) := "01111011";
			tmp(17,63) := "01111101";
			tmp(17,64) := "01111100";
			tmp(17,65) := "01111100";
			tmp(17,66) := "01111110";
			tmp(17,67) := "01101100";
			tmp(17,68) := "01110101";
			tmp(17,69) := "01111001";
			tmp(17,70) := "01110001";
			tmp(17,71) := "10000111";
			tmp(17,72) := "10010000";
			tmp(17,73) := "10001110";
			tmp(17,74) := "11000011";
			tmp(17,75) := "11101011";
			tmp(17,76) := "11111011";
			tmp(17,77) := "11111100";
			tmp(17,78) := "11111111";
			tmp(17,79) := "11111111";
			tmp(17,80) := "11111100";
			tmp(18,1) := "11111111";
			tmp(18,2) := "11111111";
			tmp(18,3) := "11111111";
			tmp(18,4) := "11111111";
			tmp(18,5) := "11111111";
			tmp(18,6) := "11111111";
			tmp(18,7) := "11111111";
			tmp(18,8) := "11111111";
			tmp(18,9) := "11111111";
			tmp(18,10) := "11111111";
			tmp(18,11) := "11111111";
			tmp(18,12) := "11111111";
			tmp(18,13) := "11111111";
			tmp(18,14) := "11111111";
			tmp(18,15) := "11111111";
			tmp(18,16) := "11111111";
			tmp(18,17) := "11111111";
			tmp(18,18) := "11111111";
			tmp(18,19) := "11111100";
			tmp(18,20) := "11111100";
			tmp(18,21) := "11111100";
			tmp(18,22) := "11111110";
			tmp(18,23) := "11111111";
			tmp(18,24) := "11111111";
			tmp(18,25) := "11110110";
			tmp(18,26) := "11111111";
			tmp(18,27) := "11111111";
			tmp(18,28) := "11111101";
			tmp(18,29) := "11111110";
			tmp(18,30) := "11111000";
			tmp(18,31) := "11110000";
			tmp(18,32) := "11011011";
			tmp(18,33) := "11011110";
			tmp(18,34) := "11010111";
			tmp(18,35) := "11010100";
			tmp(18,36) := "11001011";
			tmp(18,37) := "11001010";
			tmp(18,38) := "11001001";
			tmp(18,39) := "11010101";
			tmp(18,40) := "11000011";
			tmp(18,41) := "11000001";
			tmp(18,42) := "11000010";
			tmp(18,43) := "11001111";
			tmp(18,44) := "11010010";
			tmp(18,45) := "10111001";
			tmp(18,46) := "10101001";
			tmp(18,47) := "10011110";
			tmp(18,48) := "10100010";
			tmp(18,49) := "10011011";
			tmp(18,50) := "10010100";
			tmp(18,51) := "10100100";
			tmp(18,52) := "10101000";
			tmp(18,53) := "10011010";
			tmp(18,54) := "10001000";
			tmp(18,55) := "10001001";
			tmp(18,56) := "10001011";
			tmp(18,57) := "01111011";
			tmp(18,58) := "01111011";
			tmp(18,59) := "10000000";
			tmp(18,60) := "10000010";
			tmp(18,61) := "10000011";
			tmp(18,62) := "01111010";
			tmp(18,63) := "01111010";
			tmp(18,64) := "01111010";
			tmp(18,65) := "10000001";
			tmp(18,66) := "01111011";
			tmp(18,67) := "01101001";
			tmp(18,68) := "01101010";
			tmp(18,69) := "01100100";
			tmp(18,70) := "01101110";
			tmp(18,71) := "01110111";
			tmp(18,72) := "10000000";
			tmp(18,73) := "10001101";
			tmp(18,74) := "10100001";
			tmp(18,75) := "11010001";
			tmp(18,76) := "11111001";
			tmp(18,77) := "11111111";
			tmp(18,78) := "11111111";
			tmp(18,79) := "11111100";
			tmp(18,80) := "11111100";
			tmp(19,1) := "11111111";
			tmp(19,2) := "11111111";
			tmp(19,3) := "11111111";
			tmp(19,4) := "11111111";
			tmp(19,5) := "11111111";
			tmp(19,6) := "11111111";
			tmp(19,7) := "11111111";
			tmp(19,8) := "11111111";
			tmp(19,9) := "11111111";
			tmp(19,10) := "11111111";
			tmp(19,11) := "11111111";
			tmp(19,12) := "11111111";
			tmp(19,13) := "11111111";
			tmp(19,14) := "11111111";
			tmp(19,15) := "11111111";
			tmp(19,16) := "11111111";
			tmp(19,17) := "11111111";
			tmp(19,18) := "11111110";
			tmp(19,19) := "11111110";
			tmp(19,20) := "11111100";
			tmp(19,21) := "11111110";
			tmp(19,22) := "11111111";
			tmp(19,23) := "11111010";
			tmp(19,24) := "11111001";
			tmp(19,25) := "11111111";
			tmp(19,26) := "11111110";
			tmp(19,27) := "11111111";
			tmp(19,28) := "11111100";
			tmp(19,29) := "11110101";
			tmp(19,30) := "11101001";
			tmp(19,31) := "11101100";
			tmp(19,32) := "11011011";
			tmp(19,33) := "11010111";
			tmp(19,34) := "11010011";
			tmp(19,35) := "11010110";
			tmp(19,36) := "11010001";
			tmp(19,37) := "11001011";
			tmp(19,38) := "11010010";
			tmp(19,39) := "11000101";
			tmp(19,40) := "10111110";
			tmp(19,41) := "10111011";
			tmp(19,42) := "10110101";
			tmp(19,43) := "10110011";
			tmp(19,44) := "11000010";
			tmp(19,45) := "10101111";
			tmp(19,46) := "10001111";
			tmp(19,47) := "10001100";
			tmp(19,48) := "10010101";
			tmp(19,49) := "10001101";
			tmp(19,50) := "10000011";
			tmp(19,51) := "10000111";
			tmp(19,52) := "10100000";
			tmp(19,53) := "10010000";
			tmp(19,54) := "10000010";
			tmp(19,55) := "01111010";
			tmp(19,56) := "01111011";
			tmp(19,57) := "01111010";
			tmp(19,58) := "01110011";
			tmp(19,59) := "01110010";
			tmp(19,60) := "10000010";
			tmp(19,61) := "10000001";
			tmp(19,62) := "01110110";
			tmp(19,63) := "01110101";
			tmp(19,64) := "10000011";
			tmp(19,65) := "01111001";
			tmp(19,66) := "01101010";
			tmp(19,67) := "01100001";
			tmp(19,68) := "01100001";
			tmp(19,69) := "01101011";
			tmp(19,70) := "01100100";
			tmp(19,71) := "01111001";
			tmp(19,72) := "01111100";
			tmp(19,73) := "10000111";
			tmp(19,74) := "10010111";
			tmp(19,75) := "10101101";
			tmp(19,76) := "11101101";
			tmp(19,77) := "11111110";
			tmp(19,78) := "11111110";
			tmp(19,79) := "11111111";
			tmp(19,80) := "11111111";
			tmp(20,1) := "11111111";
			tmp(20,2) := "11111111";
			tmp(20,3) := "11111111";
			tmp(20,4) := "11111111";
			tmp(20,5) := "11111111";
			tmp(20,6) := "11111111";
			tmp(20,7) := "11111111";
			tmp(20,8) := "11111111";
			tmp(20,9) := "11111111";
			tmp(20,10) := "11111111";
			tmp(20,11) := "11111111";
			tmp(20,12) := "11111111";
			tmp(20,13) := "11111111";
			tmp(20,14) := "11111111";
			tmp(20,15) := "11111111";
			tmp(20,16) := "11111111";
			tmp(20,17) := "11111100";
			tmp(20,18) := "11111111";
			tmp(20,19) := "11111111";
			tmp(20,20) := "11111111";
			tmp(20,21) := "11111101";
			tmp(20,22) := "11111111";
			tmp(20,23) := "11111111";
			tmp(20,24) := "11111011";
			tmp(20,25) := "11111111";
			tmp(20,26) := "11111101";
			tmp(20,27) := "11110011";
			tmp(20,28) := "11101101";
			tmp(20,29) := "11101100";
			tmp(20,30) := "11100010";
			tmp(20,31) := "11100011";
			tmp(20,32) := "11011101";
			tmp(20,33) := "11001010";
			tmp(20,34) := "11010010";
			tmp(20,35) := "11001111";
			tmp(20,36) := "11010001";
			tmp(20,37) := "11010000";
			tmp(20,38) := "11000010";
			tmp(20,39) := "10111100";
			tmp(20,40) := "10111110";
			tmp(20,41) := "10110100";
			tmp(20,42) := "10110100";
			tmp(20,43) := "10111111";
			tmp(20,44) := "10111111";
			tmp(20,45) := "10101111";
			tmp(20,46) := "10001111";
			tmp(20,47) := "10010111";
			tmp(20,48) := "10010011";
			tmp(20,49) := "10010001";
			tmp(20,50) := "10000110";
			tmp(20,51) := "10000011";
			tmp(20,52) := "10001101";
			tmp(20,53) := "10000111";
			tmp(20,54) := "01110111";
			tmp(20,55) := "01111000";
			tmp(20,56) := "01110110";
			tmp(20,57) := "01110000";
			tmp(20,58) := "01110000";
			tmp(20,59) := "01101111";
			tmp(20,60) := "01110001";
			tmp(20,61) := "01111101";
			tmp(20,62) := "01110001";
			tmp(20,63) := "01101111";
			tmp(20,64) := "01101100";
			tmp(20,65) := "01110110";
			tmp(20,66) := "01101100";
			tmp(20,67) := "01101000";
			tmp(20,68) := "01101111";
			tmp(20,69) := "01111001";
			tmp(20,70) := "01111001";
			tmp(20,71) := "01111010";
			tmp(20,72) := "01111100";
			tmp(20,73) := "10010100";
			tmp(20,74) := "10010001";
			tmp(20,75) := "10000110";
			tmp(20,76) := "11011011";
			tmp(20,77) := "11111011";
			tmp(20,78) := "11111111";
			tmp(20,79) := "11111110";
			tmp(20,80) := "11111111";
			tmp(21,1) := "11111111";
			tmp(21,2) := "11111111";
			tmp(21,3) := "11111111";
			tmp(21,4) := "11111111";
			tmp(21,5) := "11111111";
			tmp(21,6) := "11111111";
			tmp(21,7) := "11111111";
			tmp(21,8) := "11111111";
			tmp(21,9) := "11111111";
			tmp(21,10) := "11111111";
			tmp(21,11) := "11111111";
			tmp(21,12) := "11111111";
			tmp(21,13) := "11111111";
			tmp(21,14) := "11111111";
			tmp(21,15) := "11111111";
			tmp(21,16) := "11111111";
			tmp(21,17) := "11111111";
			tmp(21,18) := "11111111";
			tmp(21,19) := "11111111";
			tmp(21,20) := "11111111";
			tmp(21,21) := "11111111";
			tmp(21,22) := "11111111";
			tmp(21,23) := "11111111";
			tmp(21,24) := "11111111";
			tmp(21,25) := "11111111";
			tmp(21,26) := "11111010";
			tmp(21,27) := "11110001";
			tmp(21,28) := "11100000";
			tmp(21,29) := "11011101";
			tmp(21,30) := "11011000";
			tmp(21,31) := "11011111";
			tmp(21,32) := "11000010";
			tmp(21,33) := "11010000";
			tmp(21,34) := "11001101";
			tmp(21,35) := "11001001";
			tmp(21,36) := "11001101";
			tmp(21,37) := "11010001";
			tmp(21,38) := "10111011";
			tmp(21,39) := "10111010";
			tmp(21,40) := "10110010";
			tmp(21,41) := "10101111";
			tmp(21,42) := "10110111";
			tmp(21,43) := "11001010";
			tmp(21,44) := "10111001";
			tmp(21,45) := "10011100";
			tmp(21,46) := "10001011";
			tmp(21,47) := "10010011";
			tmp(21,48) := "10010111";
			tmp(21,49) := "10001100";
			tmp(21,50) := "10010001";
			tmp(21,51) := "10001011";
			tmp(21,52) := "10001011";
			tmp(21,53) := "01111110";
			tmp(21,54) := "01111101";
			tmp(21,55) := "01110111";
			tmp(21,56) := "01110100";
			tmp(21,57) := "01101100";
			tmp(21,58) := "01110001";
			tmp(21,59) := "01101010";
			tmp(21,60) := "01110010";
			tmp(21,61) := "01110010";
			tmp(21,62) := "01110000";
			tmp(21,63) := "01110000";
			tmp(21,64) := "01110010";
			tmp(21,65) := "01101011";
			tmp(21,66) := "01100110";
			tmp(21,67) := "01100001";
			tmp(21,68) := "01110100";
			tmp(21,69) := "01111100";
			tmp(21,70) := "01110010";
			tmp(21,71) := "01110110";
			tmp(21,72) := "01110100";
			tmp(21,73) := "10001000";
			tmp(21,74) := "10001101";
			tmp(21,75) := "10001111";
			tmp(21,76) := "10111010";
			tmp(21,77) := "11111110";
			tmp(21,78) := "11111111";
			tmp(21,79) := "11111111";
			tmp(21,80) := "11111010";
			tmp(22,1) := "11111111";
			tmp(22,2) := "11111111";
			tmp(22,3) := "11111111";
			tmp(22,4) := "11111111";
			tmp(22,5) := "11111111";
			tmp(22,6) := "11111111";
			tmp(22,7) := "11111111";
			tmp(22,8) := "11111111";
			tmp(22,9) := "11111111";
			tmp(22,10) := "11111111";
			tmp(22,11) := "11111111";
			tmp(22,12) := "11111111";
			tmp(22,13) := "11111111";
			tmp(22,14) := "11111111";
			tmp(22,15) := "11111111";
			tmp(22,16) := "11111111";
			tmp(22,17) := "11111111";
			tmp(22,18) := "11111111";
			tmp(22,19) := "11111100";
			tmp(22,20) := "11111111";
			tmp(22,21) := "11111111";
			tmp(22,22) := "11111011";
			tmp(22,23) := "11111011";
			tmp(22,24) := "11111011";
			tmp(22,25) := "11111101";
			tmp(22,26) := "11101111";
			tmp(22,27) := "11101010";
			tmp(22,28) := "11101101";
			tmp(22,29) := "11101011";
			tmp(22,30) := "11100110";
			tmp(22,31) := "11011100";
			tmp(22,32) := "11001001";
			tmp(22,33) := "11000110";
			tmp(22,34) := "11010011";
			tmp(22,35) := "11000010";
			tmp(22,36) := "11000001";
			tmp(22,37) := "11000001";
			tmp(22,38) := "10111011";
			tmp(22,39) := "10110110";
			tmp(22,40) := "10101110";
			tmp(22,41) := "10100111";
			tmp(22,42) := "10100111";
			tmp(22,43) := "10101011";
			tmp(22,44) := "10100001";
			tmp(22,45) := "10010111";
			tmp(22,46) := "10001100";
			tmp(22,47) := "10010000";
			tmp(22,48) := "10010010";
			tmp(22,49) := "10000000";
			tmp(22,50) := "10000011";
			tmp(22,51) := "10000111";
			tmp(22,52) := "01111001";
			tmp(22,53) := "01110111";
			tmp(22,54) := "01101110";
			tmp(22,55) := "01101011";
			tmp(22,56) := "01100101";
			tmp(22,57) := "01100011";
			tmp(22,58) := "01100110";
			tmp(22,59) := "01101011";
			tmp(22,60) := "01100111";
			tmp(22,61) := "01101100";
			tmp(22,62) := "01100110";
			tmp(22,63) := "01110000";
			tmp(22,64) := "01110001";
			tmp(22,65) := "01101001";
			tmp(22,66) := "01101101";
			tmp(22,67) := "10000011";
			tmp(22,68) := "01111000";
			tmp(22,69) := "01110111";
			tmp(22,70) := "01110101";
			tmp(22,71) := "01111011";
			tmp(22,72) := "01111000";
			tmp(22,73) := "10000001";
			tmp(22,74) := "01111101";
			tmp(22,75) := "10000101";
			tmp(22,76) := "10101001";
			tmp(22,77) := "11100111";
			tmp(22,78) := "11111110";
			tmp(22,79) := "11111110";
			tmp(22,80) := "11111111";
			tmp(23,1) := "11111111";
			tmp(23,2) := "11111111";
			tmp(23,3) := "11111111";
			tmp(23,4) := "11111111";
			tmp(23,5) := "11111111";
			tmp(23,6) := "11111111";
			tmp(23,7) := "11111111";
			tmp(23,8) := "11111111";
			tmp(23,9) := "11111111";
			tmp(23,10) := "11111111";
			tmp(23,11) := "11111111";
			tmp(23,12) := "11111111";
			tmp(23,13) := "11111111";
			tmp(23,14) := "11111111";
			tmp(23,15) := "11111111";
			tmp(23,16) := "11111111";
			tmp(23,17) := "11111110";
			tmp(23,18) := "11111110";
			tmp(23,19) := "11111100";
			tmp(23,20) := "11111111";
			tmp(23,21) := "11111010";
			tmp(23,22) := "11111011";
			tmp(23,23) := "11111111";
			tmp(23,24) := "11101111";
			tmp(23,25) := "11101100";
			tmp(23,26) := "11101101";
			tmp(23,27) := "11101011";
			tmp(23,28) := "11100111";
			tmp(23,29) := "11011101";
			tmp(23,30) := "11100011";
			tmp(23,31) := "11011011";
			tmp(23,32) := "11010101";
			tmp(23,33) := "11001100";
			tmp(23,34) := "11010001";
			tmp(23,35) := "11001101";
			tmp(23,36) := "10111101";
			tmp(23,37) := "10101100";
			tmp(23,38) := "10111111";
			tmp(23,39) := "10111010";
			tmp(23,40) := "10101010";
			tmp(23,41) := "10011011";
			tmp(23,42) := "10010011";
			tmp(23,43) := "10100001";
			tmp(23,44) := "10101010";
			tmp(23,45) := "10001110";
			tmp(23,46) := "10001001";
			tmp(23,47) := "10001110";
			tmp(23,48) := "10001010";
			tmp(23,49) := "01110111";
			tmp(23,50) := "01110101";
			tmp(23,51) := "01110100";
			tmp(23,52) := "01110101";
			tmp(23,53) := "01110001";
			tmp(23,54) := "01110001";
			tmp(23,55) := "01101011";
			tmp(23,56) := "01100111";
			tmp(23,57) := "01101001";
			tmp(23,58) := "01100010";
			tmp(23,59) := "01011011";
			tmp(23,60) := "01011111";
			tmp(23,61) := "01100000";
			tmp(23,62) := "01011010";
			tmp(23,63) := "01011011";
			tmp(23,64) := "01100010";
			tmp(23,65) := "01100001";
			tmp(23,66) := "01110110";
			tmp(23,67) := "10000011";
			tmp(23,68) := "10000101";
			tmp(23,69) := "01110011";
			tmp(23,70) := "01110111";
			tmp(23,71) := "01111110";
			tmp(23,72) := "10000100";
			tmp(23,73) := "10000011";
			tmp(23,74) := "01111111";
			tmp(23,75) := "10000011";
			tmp(23,76) := "10011100";
			tmp(23,77) := "11111010";
			tmp(23,78) := "11111111";
			tmp(23,79) := "11111101";
			tmp(23,80) := "11111111";
			tmp(24,1) := "11111111";
			tmp(24,2) := "11111111";
			tmp(24,3) := "11111111";
			tmp(24,4) := "11111111";
			tmp(24,5) := "11111111";
			tmp(24,6) := "11111111";
			tmp(24,7) := "11111111";
			tmp(24,8) := "11111111";
			tmp(24,9) := "11111111";
			tmp(24,10) := "11111111";
			tmp(24,11) := "11111111";
			tmp(24,12) := "11111111";
			tmp(24,13) := "11111111";
			tmp(24,14) := "11111111";
			tmp(24,15) := "11111111";
			tmp(24,16) := "11111111";
			tmp(24,17) := "11111111";
			tmp(24,18) := "11111110";
			tmp(24,19) := "11111111";
			tmp(24,20) := "11111101";
			tmp(24,21) := "11111001";
			tmp(24,22) := "11111110";
			tmp(24,23) := "11110010";
			tmp(24,24) := "11101111";
			tmp(24,25) := "11101100";
			tmp(24,26) := "11100100";
			tmp(24,27) := "11010010";
			tmp(24,28) := "11011011";
			tmp(24,29) := "11100001";
			tmp(24,30) := "11001100";
			tmp(24,31) := "11000110";
			tmp(24,32) := "11000111";
			tmp(24,33) := "11011001";
			tmp(24,34) := "11010110";
			tmp(24,35) := "11001111";
			tmp(24,36) := "11000101";
			tmp(24,37) := "10110110";
			tmp(24,38) := "10111101";
			tmp(24,39) := "10111010";
			tmp(24,40) := "10110001";
			tmp(24,41) := "10011101";
			tmp(24,42) := "10010110";
			tmp(24,43) := "10011110";
			tmp(24,44) := "10010110";
			tmp(24,45) := "10000101";
			tmp(24,46) := "10001110";
			tmp(24,47) := "10001011";
			tmp(24,48) := "10001001";
			tmp(24,49) := "01111111";
			tmp(24,50) := "01111001";
			tmp(24,51) := "01110110";
			tmp(24,52) := "01110010";
			tmp(24,53) := "01101011";
			tmp(24,54) := "01101101";
			tmp(24,55) := "01101010";
			tmp(24,56) := "01100110";
			tmp(24,57) := "01100010";
			tmp(24,58) := "01100101";
			tmp(24,59) := "01100001";
			tmp(24,60) := "01011011";
			tmp(24,61) := "01011111";
			tmp(24,62) := "01011111";
			tmp(24,63) := "01100010";
			tmp(24,64) := "01100100";
			tmp(24,65) := "01100111";
			tmp(24,66) := "01110111";
			tmp(24,67) := "01111011";
			tmp(24,68) := "01110110";
			tmp(24,69) := "01110001";
			tmp(24,70) := "01101110";
			tmp(24,71) := "01110010";
			tmp(24,72) := "01101101";
			tmp(24,73) := "01111111";
			tmp(24,74) := "01111101";
			tmp(24,75) := "10001001";
			tmp(24,76) := "10110001";
			tmp(24,77) := "11100010";
			tmp(24,78) := "11111111";
			tmp(24,79) := "11111100";
			tmp(24,80) := "11111111";
			tmp(25,1) := "11111111";
			tmp(25,2) := "11111111";
			tmp(25,3) := "11111111";
			tmp(25,4) := "11111111";
			tmp(25,5) := "11111111";
			tmp(25,6) := "11111111";
			tmp(25,7) := "11111111";
			tmp(25,8) := "11111111";
			tmp(25,9) := "11111111";
			tmp(25,10) := "11111101";
			tmp(25,11) := "11111100";
			tmp(25,12) := "11111111";
			tmp(25,13) := "11111111";
			tmp(25,14) := "11111110";
			tmp(25,15) := "11111100";
			tmp(25,16) := "11111111";
			tmp(25,17) := "11111111";
			tmp(25,18) := "11111010";
			tmp(25,19) := "11111111";
			tmp(25,20) := "11111011";
			tmp(25,21) := "11111100";
			tmp(25,22) := "11111000";
			tmp(25,23) := "11110110";
			tmp(25,24) := "11100011";
			tmp(25,25) := "11100101";
			tmp(25,26) := "11011011";
			tmp(25,27) := "11011010";
			tmp(25,28) := "11001101";
			tmp(25,29) := "11000110";
			tmp(25,30) := "11000011";
			tmp(25,31) := "11000011";
			tmp(25,32) := "10111101";
			tmp(25,33) := "11000010";
			tmp(25,34) := "11000100";
			tmp(25,35) := "10111111";
			tmp(25,36) := "10111010";
			tmp(25,37) := "10111001";
			tmp(25,38) := "10101010";
			tmp(25,39) := "10101101";
			tmp(25,40) := "10101011";
			tmp(25,41) := "10011001";
			tmp(25,42) := "10000100";
			tmp(25,43) := "10000000";
			tmp(25,44) := "10001000";
			tmp(25,45) := "10000110";
			tmp(25,46) := "10000001";
			tmp(25,47) := "10000101";
			tmp(25,48) := "10000010";
			tmp(25,49) := "01110001";
			tmp(25,50) := "01101010";
			tmp(25,51) := "01110101";
			tmp(25,52) := "01110001";
			tmp(25,53) := "01101100";
			tmp(25,54) := "01110010";
			tmp(25,55) := "01101001";
			tmp(25,56) := "01011110";
			tmp(25,57) := "01011101";
			tmp(25,58) := "01100100";
			tmp(25,59) := "01011011";
			tmp(25,60) := "01011010";
			tmp(25,61) := "01100001";
			tmp(25,62) := "01011100";
			tmp(25,63) := "01100000";
			tmp(25,64) := "01110001";
			tmp(25,65) := "01101001";
			tmp(25,66) := "01110011";
			tmp(25,67) := "01110111";
			tmp(25,68) := "01110100";
			tmp(25,69) := "01101101";
			tmp(25,70) := "01101100";
			tmp(25,71) := "01110000";
			tmp(25,72) := "01111110";
			tmp(25,73) := "01111111";
			tmp(25,74) := "01110111";
			tmp(25,75) := "01111010";
			tmp(25,76) := "10011001";
			tmp(25,77) := "11101010";
			tmp(25,78) := "11111001";
			tmp(25,79) := "11111000";
			tmp(25,80) := "11111111";
			tmp(26,1) := "11111111";
			tmp(26,2) := "11111111";
			tmp(26,3) := "11111111";
			tmp(26,4) := "11111111";
			tmp(26,5) := "11111111";
			tmp(26,6) := "11111111";
			tmp(26,7) := "11111111";
			tmp(26,8) := "11111111";
			tmp(26,9) := "11111100";
			tmp(26,10) := "11111111";
			tmp(26,11) := "11111111";
			tmp(26,12) := "11111111";
			tmp(26,13) := "11111111";
			tmp(26,14) := "11111011";
			tmp(26,15) := "11111110";
			tmp(26,16) := "11111111";
			tmp(26,17) := "11111101";
			tmp(26,18) := "11111100";
			tmp(26,19) := "11111111";
			tmp(26,20) := "11111101";
			tmp(26,21) := "11110011";
			tmp(26,22) := "11111101";
			tmp(26,23) := "11101100";
			tmp(26,24) := "11101000";
			tmp(26,25) := "11100110";
			tmp(26,26) := "11101001";
			tmp(26,27) := "11011010";
			tmp(26,28) := "11010111";
			tmp(26,29) := "11001111";
			tmp(26,30) := "11001001";
			tmp(26,31) := "11000101";
			tmp(26,32) := "11000100";
			tmp(26,33) := "11001001";
			tmp(26,34) := "10111100";
			tmp(26,35) := "11000111";
			tmp(26,36) := "10110100";
			tmp(26,37) := "10101110";
			tmp(26,38) := "10101011";
			tmp(26,39) := "10101010";
			tmp(26,40) := "10101000";
			tmp(26,41) := "10010111";
			tmp(26,42) := "10000101";
			tmp(26,43) := "10000100";
			tmp(26,44) := "10000100";
			tmp(26,45) := "01111001";
			tmp(26,46) := "01111000";
			tmp(26,47) := "10000010";
			tmp(26,48) := "10000010";
			tmp(26,49) := "01110010";
			tmp(26,50) := "01110000";
			tmp(26,51) := "01101110";
			tmp(26,52) := "01100111";
			tmp(26,53) := "01100100";
			tmp(26,54) := "01101011";
			tmp(26,55) := "01100101";
			tmp(26,56) := "01100001";
			tmp(26,57) := "01011010";
			tmp(26,58) := "01011000";
			tmp(26,59) := "01011101";
			tmp(26,60) := "01010110";
			tmp(26,61) := "01010010";
			tmp(26,62) := "01011101";
			tmp(26,63) := "01100100";
			tmp(26,64) := "01100111";
			tmp(26,65) := "01100110";
			tmp(26,66) := "01100010";
			tmp(26,67) := "01100111";
			tmp(26,68) := "01110000";
			tmp(26,69) := "01110010";
			tmp(26,70) := "01110000";
			tmp(26,71) := "01110101";
			tmp(26,72) := "10001100";
			tmp(26,73) := "10001111";
			tmp(26,74) := "10001001";
			tmp(26,75) := "10001010";
			tmp(26,76) := "10001101";
			tmp(26,77) := "10111100";
			tmp(26,78) := "11111111";
			tmp(26,79) := "11111110";
			tmp(26,80) := "11111110";
			tmp(27,1) := "11111111";
			tmp(27,2) := "11111111";
			tmp(27,3) := "11111111";
			tmp(27,4) := "11111111";
			tmp(27,5) := "11111111";
			tmp(27,6) := "11111111";
			tmp(27,7) := "11111111";
			tmp(27,8) := "11111111";
			tmp(27,9) := "11111110";
			tmp(27,10) := "11110010";
			tmp(27,11) := "11111011";
			tmp(27,12) := "11111110";
			tmp(27,13) := "11111101";
			tmp(27,14) := "11111111";
			tmp(27,15) := "11111111";
			tmp(27,16) := "11111100";
			tmp(27,17) := "11111111";
			tmp(27,18) := "11111110";
			tmp(27,19) := "11111111";
			tmp(27,20) := "11111101";
			tmp(27,21) := "11110100";
			tmp(27,22) := "11110000";
			tmp(27,23) := "11101100";
			tmp(27,24) := "11100010";
			tmp(27,25) := "11100010";
			tmp(27,26) := "11011011";
			tmp(27,27) := "11001000";
			tmp(27,28) := "11000010";
			tmp(27,29) := "11010001";
			tmp(27,30) := "11010111";
			tmp(27,31) := "11010001";
			tmp(27,32) := "11001100";
			tmp(27,33) := "11001010";
			tmp(27,34) := "11001000";
			tmp(27,35) := "10111101";
			tmp(27,36) := "10111011";
			tmp(27,37) := "10110100";
			tmp(27,38) := "10110010";
			tmp(27,39) := "10100100";
			tmp(27,40) := "10011011";
			tmp(27,41) := "10010011";
			tmp(27,42) := "10000111";
			tmp(27,43) := "10001000";
			tmp(27,44) := "10001000";
			tmp(27,45) := "01111011";
			tmp(27,46) := "01110010";
			tmp(27,47) := "01111000";
			tmp(27,48) := "01111011";
			tmp(27,49) := "01101100";
			tmp(27,50) := "01101001";
			tmp(27,51) := "01100111";
			tmp(27,52) := "01100110";
			tmp(27,53) := "01100101";
			tmp(27,54) := "01100100";
			tmp(27,55) := "01011110";
			tmp(27,56) := "01100010";
			tmp(27,57) := "01100011";
			tmp(27,58) := "01011100";
			tmp(27,59) := "01100101";
			tmp(27,60) := "01011101";
			tmp(27,61) := "01010110";
			tmp(27,62) := "01100011";
			tmp(27,63) := "01100101";
			tmp(27,64) := "01100001";
			tmp(27,65) := "01100100";
			tmp(27,66) := "01011110";
			tmp(27,67) := "01100100";
			tmp(27,68) := "01101100";
			tmp(27,69) := "01101100";
			tmp(27,70) := "01101111";
			tmp(27,71) := "01111011";
			tmp(27,72) := "10010000";
			tmp(27,73) := "10011010";
			tmp(27,74) := "10001111";
			tmp(27,75) := "10010101";
			tmp(27,76) := "10001100";
			tmp(27,77) := "10101101";
			tmp(27,78) := "11101111";
			tmp(27,79) := "11111111";
			tmp(27,80) := "11111111";
			tmp(28,1) := "11111111";
			tmp(28,2) := "11111111";
			tmp(28,3) := "11111111";
			tmp(28,4) := "11111111";
			tmp(28,5) := "11111111";
			tmp(28,6) := "11111111";
			tmp(28,7) := "11111111";
			tmp(28,8) := "11111111";
			tmp(28,9) := "11111111";
			tmp(28,10) := "11100111";
			tmp(28,11) := "10110100";
			tmp(28,12) := "11000010";
			tmp(28,13) := "11111100";
			tmp(28,14) := "11111111";
			tmp(28,15) := "11111111";
			tmp(28,16) := "11111010";
			tmp(28,17) := "11111111";
			tmp(28,18) := "11111110";
			tmp(28,19) := "11111011";
			tmp(28,20) := "11101110";
			tmp(28,21) := "11110011";
			tmp(28,22) := "11011111";
			tmp(28,23) := "11010110";
			tmp(28,24) := "11010110";
			tmp(28,25) := "11011110";
			tmp(28,26) := "11010011";
			tmp(28,27) := "11001011";
			tmp(28,28) := "11001011";
			tmp(28,29) := "11010000";
			tmp(28,30) := "11001010";
			tmp(28,31) := "11000110";
			tmp(28,32) := "11001100";
			tmp(28,33) := "11001101";
			tmp(28,34) := "10110111";
			tmp(28,35) := "10110111";
			tmp(28,36) := "10100101";
			tmp(28,37) := "10100110";
			tmp(28,38) := "10100000";
			tmp(28,39) := "10010111";
			tmp(28,40) := "10010101";
			tmp(28,41) := "10001001";
			tmp(28,42) := "01111000";
			tmp(28,43) := "01111111";
			tmp(28,44) := "10000101";
			tmp(28,45) := "01110110";
			tmp(28,46) := "01110011";
			tmp(28,47) := "01111011";
			tmp(28,48) := "01110101";
			tmp(28,49) := "01100111";
			tmp(28,50) := "01100110";
			tmp(28,51) := "01101010";
			tmp(28,52) := "01100110";
			tmp(28,53) := "01100000";
			tmp(28,54) := "01100000";
			tmp(28,55) := "01100000";
			tmp(28,56) := "01101010";
			tmp(28,57) := "01101011";
			tmp(28,58) := "01100110";
			tmp(28,59) := "01100010";
			tmp(28,60) := "01011100";
			tmp(28,61) := "01011010";
			tmp(28,62) := "01011111";
			tmp(28,63) := "01011111";
			tmp(28,64) := "01010111";
			tmp(28,65) := "01011000";
			tmp(28,66) := "01011000";
			tmp(28,67) := "01101001";
			tmp(28,68) := "01111100";
			tmp(28,69) := "10000001";
			tmp(28,70) := "10000101";
			tmp(28,71) := "10001111";
			tmp(28,72) := "10011010";
			tmp(28,73) := "10001000";
			tmp(28,74) := "10001000";
			tmp(28,75) := "10010000";
			tmp(28,76) := "10001010";
			tmp(28,77) := "10010001";
			tmp(28,78) := "11001101";
			tmp(28,79) := "11111111";
			tmp(28,80) := "11111100";
			tmp(29,1) := "11111111";
			tmp(29,2) := "11111111";
			tmp(29,3) := "11111111";
			tmp(29,4) := "11111111";
			tmp(29,5) := "11111111";
			tmp(29,6) := "11111111";
			tmp(29,7) := "11111111";
			tmp(29,8) := "11111111";
			tmp(29,9) := "11111111";
			tmp(29,10) := "11111111";
			tmp(29,11) := "11011111";
			tmp(29,12) := "10001001";
			tmp(29,13) := "11000110";
			tmp(29,14) := "11111100";
			tmp(29,15) := "11111111";
			tmp(29,16) := "11111110";
			tmp(29,17) := "11111111";
			tmp(29,18) := "11111111";
			tmp(29,19) := "11111001";
			tmp(29,20) := "11111011";
			tmp(29,21) := "11110101";
			tmp(29,22) := "11100101";
			tmp(29,23) := "11011011";
			tmp(29,24) := "11011010";
			tmp(29,25) := "11011010";
			tmp(29,26) := "11010111";
			tmp(29,27) := "11001011";
			tmp(29,28) := "11000101";
			tmp(29,29) := "11010100";
			tmp(29,30) := "11000011";
			tmp(29,31) := "11000101";
			tmp(29,32) := "11000010";
			tmp(29,33) := "10111011";
			tmp(29,34) := "11000000";
			tmp(29,35) := "10110011";
			tmp(29,36) := "10100011";
			tmp(29,37) := "10011110";
			tmp(29,38) := "10010100";
			tmp(29,39) := "10011000";
			tmp(29,40) := "10010010";
			tmp(29,41) := "10000001";
			tmp(29,42) := "01111001";
			tmp(29,43) := "01111011";
			tmp(29,44) := "01111010";
			tmp(29,45) := "01111010";
			tmp(29,46) := "01110101";
			tmp(29,47) := "01110001";
			tmp(29,48) := "01100111";
			tmp(29,49) := "01100101";
			tmp(29,50) := "01101010";
			tmp(29,51) := "01101010";
			tmp(29,52) := "01100101";
			tmp(29,53) := "01100100";
			tmp(29,54) := "01101001";
			tmp(29,55) := "01101010";
			tmp(29,56) := "01101011";
			tmp(29,57) := "01011010";
			tmp(29,58) := "01011101";
			tmp(29,59) := "01011001";
			tmp(29,60) := "01011010";
			tmp(29,61) := "01011101";
			tmp(29,62) := "01100010";
			tmp(29,63) := "01100011";
			tmp(29,64) := "01010111";
			tmp(29,65) := "01011010";
			tmp(29,66) := "01101100";
			tmp(29,67) := "01110100";
			tmp(29,68) := "10000100";
			tmp(29,69) := "10010101";
			tmp(29,70) := "10011011";
			tmp(29,71) := "10100010";
			tmp(29,72) := "10100001";
			tmp(29,73) := "10001101";
			tmp(29,74) := "10000011";
			tmp(29,75) := "10001111";
			tmp(29,76) := "10001100";
			tmp(29,77) := "10010101";
			tmp(29,78) := "10110011";
			tmp(29,79) := "11110000";
			tmp(29,80) := "11111010";
			tmp(30,1) := "11111111";
			tmp(30,2) := "11111111";
			tmp(30,3) := "11111111";
			tmp(30,4) := "11111111";
			tmp(30,5) := "11111111";
			tmp(30,6) := "11111111";
			tmp(30,7) := "11111111";
			tmp(30,8) := "11111111";
			tmp(30,9) := "11111110";
			tmp(30,10) := "11111111";
			tmp(30,11) := "11111000";
			tmp(30,12) := "11100011";
			tmp(30,13) := "01110001";
			tmp(30,14) := "10110110";
			tmp(30,15) := "11111001";
			tmp(30,16) := "11111111";
			tmp(30,17) := "11111011";
			tmp(30,18) := "11111111";
			tmp(30,19) := "11110110";
			tmp(30,20) := "11110111";
			tmp(30,21) := "11110100";
			tmp(30,22) := "11100111";
			tmp(30,23) := "11100000";
			tmp(30,24) := "11010111";
			tmp(30,25) := "11011100";
			tmp(30,26) := "11100101";
			tmp(30,27) := "11001110";
			tmp(30,28) := "11001010";
			tmp(30,29) := "11000011";
			tmp(30,30) := "11010001";
			tmp(30,31) := "11001100";
			tmp(30,32) := "11000111";
			tmp(30,33) := "10111101";
			tmp(30,34) := "11001001";
			tmp(30,35) := "10111100";
			tmp(30,36) := "10101111";
			tmp(30,37) := "10101010";
			tmp(30,38) := "10010111";
			tmp(30,39) := "10010100";
			tmp(30,40) := "10010000";
			tmp(30,41) := "10001100";
			tmp(30,42) := "10000010";
			tmp(30,43) := "10000000";
			tmp(30,44) := "01111111";
			tmp(30,45) := "01111011";
			tmp(30,46) := "01110110";
			tmp(30,47) := "01101101";
			tmp(30,48) := "01100010";
			tmp(30,49) := "01100101";
			tmp(30,50) := "01101011";
			tmp(30,51) := "01100011";
			tmp(30,52) := "01100010";
			tmp(30,53) := "01100100";
			tmp(30,54) := "01100100";
			tmp(30,55) := "01100110";
			tmp(30,56) := "01100001";
			tmp(30,57) := "01010011";
			tmp(30,58) := "01010111";
			tmp(30,59) := "01010110";
			tmp(30,60) := "01010110";
			tmp(30,61) := "01011111";
			tmp(30,62) := "01100100";
			tmp(30,63) := "01100011";
			tmp(30,64) := "01100111";
			tmp(30,65) := "01100001";
			tmp(30,66) := "01110110";
			tmp(30,67) := "10000100";
			tmp(30,68) := "10001010";
			tmp(30,69) := "10001100";
			tmp(30,70) := "10011011";
			tmp(30,71) := "10101001";
			tmp(30,72) := "10010101";
			tmp(30,73) := "10010001";
			tmp(30,74) := "10010101";
			tmp(30,75) := "10010101";
			tmp(30,76) := "10010111";
			tmp(30,77) := "10010110";
			tmp(30,78) := "10100000";
			tmp(30,79) := "11110011";
			tmp(30,80) := "11111111";
			tmp(31,1) := "11111111";
			tmp(31,2) := "11111111";
			tmp(31,3) := "11111111";
			tmp(31,4) := "11111111";
			tmp(31,5) := "11111111";
			tmp(31,6) := "11111111";
			tmp(31,7) := "11111111";
			tmp(31,8) := "11111111";
			tmp(31,9) := "11111100";
			tmp(31,10) := "11111111";
			tmp(31,11) := "11111111";
			tmp(31,12) := "11111110";
			tmp(31,13) := "11000000";
			tmp(31,14) := "01100011";
			tmp(31,15) := "10110101";
			tmp(31,16) := "11111000";
			tmp(31,17) := "11111111";
			tmp(31,18) := "11110001";
			tmp(31,19) := "11111000";
			tmp(31,20) := "11110111";
			tmp(31,21) := "11101100";
			tmp(31,22) := "11100001";
			tmp(31,23) := "11100010";
			tmp(31,24) := "11100100";
			tmp(31,25) := "11101011";
			tmp(31,26) := "11100010";
			tmp(31,27) := "11010110";
			tmp(31,28) := "11010010";
			tmp(31,29) := "11000100";
			tmp(31,30) := "11000011";
			tmp(31,31) := "10111110";
			tmp(31,32) := "10110110";
			tmp(31,33) := "10110011";
			tmp(31,34) := "10110110";
			tmp(31,35) := "10101111";
			tmp(31,36) := "10101110";
			tmp(31,37) := "10011011";
			tmp(31,38) := "10011111";
			tmp(31,39) := "10010101";
			tmp(31,40) := "10001001";
			tmp(31,41) := "10001010";
			tmp(31,42) := "10000110";
			tmp(31,43) := "10000011";
			tmp(31,44) := "10000000";
			tmp(31,45) := "01111110";
			tmp(31,46) := "01110011";
			tmp(31,47) := "01100110";
			tmp(31,48) := "01100001";
			tmp(31,49) := "01100011";
			tmp(31,50) := "01100100";
			tmp(31,51) := "01100011";
			tmp(31,52) := "01100100";
			tmp(31,53) := "01100001";
			tmp(31,54) := "01100000";
			tmp(31,55) := "01100010";
			tmp(31,56) := "01100100";
			tmp(31,57) := "01011001";
			tmp(31,58) := "01010111";
			tmp(31,59) := "01011000";
			tmp(31,60) := "01011100";
			tmp(31,61) := "01011111";
			tmp(31,62) := "01011100";
			tmp(31,63) := "01011100";
			tmp(31,64) := "01101010";
			tmp(31,65) := "01111101";
			tmp(31,66) := "10010000";
			tmp(31,67) := "10001110";
			tmp(31,68) := "10001011";
			tmp(31,69) := "10010000";
			tmp(31,70) := "10001110";
			tmp(31,71) := "10010011";
			tmp(31,72) := "10001100";
			tmp(31,73) := "10000110";
			tmp(31,74) := "10010011";
			tmp(31,75) := "10001010";
			tmp(31,76) := "10000011";
			tmp(31,77) := "10001111";
			tmp(31,78) := "10011111";
			tmp(31,79) := "11011010";
			tmp(31,80) := "11111100";
			tmp(32,1) := "11111111";
			tmp(32,2) := "11111111";
			tmp(32,3) := "11111111";
			tmp(32,4) := "11111111";
			tmp(32,5) := "11111111";
			tmp(32,6) := "11111111";
			tmp(32,7) := "11111111";
			tmp(32,8) := "11111111";
			tmp(32,9) := "11111111";
			tmp(32,10) := "11111111";
			tmp(32,11) := "11111111";
			tmp(32,12) := "11111111";
			tmp(32,13) := "11101100";
			tmp(32,14) := "01111010";
			tmp(32,15) := "01011110";
			tmp(32,16) := "11000011";
			tmp(32,17) := "11111101";
			tmp(32,18) := "11111110";
			tmp(32,19) := "11101110";
			tmp(32,20) := "11101100";
			tmp(32,21) := "11101100";
			tmp(32,22) := "11100001";
			tmp(32,23) := "11010011";
			tmp(32,24) := "11100001";
			tmp(32,25) := "11101010";
			tmp(32,26) := "11100011";
			tmp(32,27) := "11001001";
			tmp(32,28) := "11010010";
			tmp(32,29) := "11010000";
			tmp(32,30) := "11000100";
			tmp(32,31) := "10111000";
			tmp(32,32) := "10110000";
			tmp(32,33) := "10110111";
			tmp(32,34) := "10110100";
			tmp(32,35) := "10110011";
			tmp(32,36) := "10011101";
			tmp(32,37) := "10010011";
			tmp(32,38) := "10010011";
			tmp(32,39) := "10011011";
			tmp(32,40) := "10001101";
			tmp(32,41) := "10000100";
			tmp(32,42) := "10000000";
			tmp(32,43) := "01111111";
			tmp(32,44) := "01110111";
			tmp(32,45) := "01101101";
			tmp(32,46) := "01101010";
			tmp(32,47) := "01101001";
			tmp(32,48) := "01100010";
			tmp(32,49) := "01100010";
			tmp(32,50) := "01011100";
			tmp(32,51) := "01101010";
			tmp(32,52) := "01101011";
			tmp(32,53) := "01100111";
			tmp(32,54) := "01101011";
			tmp(32,55) := "01100000";
			tmp(32,56) := "01011001";
			tmp(32,57) := "01010111";
			tmp(32,58) := "01001100";
			tmp(32,59) := "01010011";
			tmp(32,60) := "01011110";
			tmp(32,61) := "01011001";
			tmp(32,62) := "01011000";
			tmp(32,63) := "01101011";
			tmp(32,64) := "01110100";
			tmp(32,65) := "10001000";
			tmp(32,66) := "10001010";
			tmp(32,67) := "10000111";
			tmp(32,68) := "10000110";
			tmp(32,69) := "10001010";
			tmp(32,70) := "10010000";
			tmp(32,71) := "10010101";
			tmp(32,72) := "10000010";
			tmp(32,73) := "10000110";
			tmp(32,74) := "10001110";
			tmp(32,75) := "10000110";
			tmp(32,76) := "01111101";
			tmp(32,77) := "10000011";
			tmp(32,78) := "10010100";
			tmp(32,79) := "11101011";
			tmp(32,80) := "11111101";
			tmp(33,1) := "11111111";
			tmp(33,2) := "11111111";
			tmp(33,3) := "11111111";
			tmp(33,4) := "11111111";
			tmp(33,5) := "11111111";
			tmp(33,6) := "11111111";
			tmp(33,7) := "11111111";
			tmp(33,8) := "11111111";
			tmp(33,9) := "11111111";
			tmp(33,10) := "11111000";
			tmp(33,11) := "11111011";
			tmp(33,12) := "11111111";
			tmp(33,13) := "11100111";
			tmp(33,14) := "01111011";
			tmp(33,15) := "01010111";
			tmp(33,16) := "10000010";
			tmp(33,17) := "11100000";
			tmp(33,18) := "11111100";
			tmp(33,19) := "11110011";
			tmp(33,20) := "11101110";
			tmp(33,21) := "11101111";
			tmp(33,22) := "11010101";
			tmp(33,23) := "11010110";
			tmp(33,24) := "11011000";
			tmp(33,25) := "11010110";
			tmp(33,26) := "11010001";
			tmp(33,27) := "11001000";
			tmp(33,28) := "11010100";
			tmp(33,29) := "11010011";
			tmp(33,30) := "11001100";
			tmp(33,31) := "10111011";
			tmp(33,32) := "10111011";
			tmp(33,33) := "11000110";
			tmp(33,34) := "10111101";
			tmp(33,35) := "10100010";
			tmp(33,36) := "10011001";
			tmp(33,37) := "10010101";
			tmp(33,38) := "10010110";
			tmp(33,39) := "10010101";
			tmp(33,40) := "10000110";
			tmp(33,41) := "01111110";
			tmp(33,42) := "10000001";
			tmp(33,43) := "01111010";
			tmp(33,44) := "01110000";
			tmp(33,45) := "01100111";
			tmp(33,46) := "01101000";
			tmp(33,47) := "01101010";
			tmp(33,48) := "01101010";
			tmp(33,49) := "01100110";
			tmp(33,50) := "01101000";
			tmp(33,51) := "01101101";
			tmp(33,52) := "01101010";
			tmp(33,53) := "01101000";
			tmp(33,54) := "01101101";
			tmp(33,55) := "01100110";
			tmp(33,56) := "01010010";
			tmp(33,57) := "01001011";
			tmp(33,58) := "01001100";
			tmp(33,59) := "01011001";
			tmp(33,60) := "01100000";
			tmp(33,61) := "01100011";
			tmp(33,62) := "01110000";
			tmp(33,63) := "01111100";
			tmp(33,64) := "10001101";
			tmp(33,65) := "10001010";
			tmp(33,66) := "10001101";
			tmp(33,67) := "10000101";
			tmp(33,68) := "10000100";
			tmp(33,69) := "10001011";
			tmp(33,70) := "10001010";
			tmp(33,71) := "10010001";
			tmp(33,72) := "10010101";
			tmp(33,73) := "10001111";
			tmp(33,74) := "10001100";
			tmp(33,75) := "10010000";
			tmp(33,76) := "10001111";
			tmp(33,77) := "10001101";
			tmp(33,78) := "10011001";
			tmp(33,79) := "11010110";
			tmp(33,80) := "11111111";
			tmp(34,1) := "11111111";
			tmp(34,2) := "11111111";
			tmp(34,3) := "11111111";
			tmp(34,4) := "11111111";
			tmp(34,5) := "11111111";
			tmp(34,6) := "11111111";
			tmp(34,7) := "11111111";
			tmp(34,8) := "11111111";
			tmp(34,9) := "11111111";
			tmp(34,10) := "11111111";
			tmp(34,11) := "11111110";
			tmp(34,12) := "11111101";
			tmp(34,13) := "11111111";
			tmp(34,14) := "10100101";
			tmp(34,15) := "01001110";
			tmp(34,16) := "10100001";
			tmp(34,17) := "11111111";
			tmp(34,18) := "11111000";
			tmp(34,19) := "11110100";
			tmp(34,20) := "11100111";
			tmp(34,21) := "11101101";
			tmp(34,22) := "11100000";
			tmp(34,23) := "11010100";
			tmp(34,24) := "11010111";
			tmp(34,25) := "11010111";
			tmp(34,26) := "11010001";
			tmp(34,27) := "11010101";
			tmp(34,28) := "11010111";
			tmp(34,29) := "11010110";
			tmp(34,30) := "11010001";
			tmp(34,31) := "11001001";
			tmp(34,32) := "11000001";
			tmp(34,33) := "11001011";
			tmp(34,34) := "10110101";
			tmp(34,35) := "10100111";
			tmp(34,36) := "10100000";
			tmp(34,37) := "10011010";
			tmp(34,38) := "10010111";
			tmp(34,39) := "10001011";
			tmp(34,40) := "10000011";
			tmp(34,41) := "01111010";
			tmp(34,42) := "01110111";
			tmp(34,43) := "01110001";
			tmp(34,44) := "01101011";
			tmp(34,45) := "01101011";
			tmp(34,46) := "01101101";
			tmp(34,47) := "01101000";
			tmp(34,48) := "01100001";
			tmp(34,49) := "01100101";
			tmp(34,50) := "01101001";
			tmp(34,51) := "01110001";
			tmp(34,52) := "01100111";
			tmp(34,53) := "01011010";
			tmp(34,54) := "01011101";
			tmp(34,55) := "01010110";
			tmp(34,56) := "01001011";
			tmp(34,57) := "01001110";
			tmp(34,58) := "01010000";
			tmp(34,59) := "01010000";
			tmp(34,60) := "01100110";
			tmp(34,61) := "01110101";
			tmp(34,62) := "01111010";
			tmp(34,63) := "10000101";
			tmp(34,64) := "10000111";
			tmp(34,65) := "10001111";
			tmp(34,66) := "10001001";
			tmp(34,67) := "10001000";
			tmp(34,68) := "10001011";
			tmp(34,69) := "01111110";
			tmp(34,70) := "01111010";
			tmp(34,71) := "10001100";
			tmp(34,72) := "10001000";
			tmp(34,73) := "10000001";
			tmp(34,74) := "10000001";
			tmp(34,75) := "01111111";
			tmp(34,76) := "10001001";
			tmp(34,77) := "10001110";
			tmp(34,78) := "10010100";
			tmp(34,79) := "11101110";
			tmp(34,80) := "11111100";
			tmp(35,1) := "11111111";
			tmp(35,2) := "11111111";
			tmp(35,3) := "11111111";
			tmp(35,4) := "11111111";
			tmp(35,5) := "11111111";
			tmp(35,6) := "11111111";
			tmp(35,7) := "11111111";
			tmp(35,8) := "11111111";
			tmp(35,9) := "11111100";
			tmp(35,10) := "11111101";
			tmp(35,11) := "11111110";
			tmp(35,12) := "11111100";
			tmp(35,13) := "11111111";
			tmp(35,14) := "11100001";
			tmp(35,15) := "01010000";
			tmp(35,16) := "10111110";
			tmp(35,17) := "11110110";
			tmp(35,18) := "11110001";
			tmp(35,19) := "11110001";
			tmp(35,20) := "11101010";
			tmp(35,21) := "11110100";
			tmp(35,22) := "11100101";
			tmp(35,23) := "11011001";
			tmp(35,24) := "11011010";
			tmp(35,25) := "11100001";
			tmp(35,26) := "11010101";
			tmp(35,27) := "11010010";
			tmp(35,28) := "11100110";
			tmp(35,29) := "11100000";
			tmp(35,30) := "11000111";
			tmp(35,31) := "10111000";
			tmp(35,32) := "11001000";
			tmp(35,33) := "10111101";
			tmp(35,34) := "10101100";
			tmp(35,35) := "10100111";
			tmp(35,36) := "10100001";
			tmp(35,37) := "10010100";
			tmp(35,38) := "10000110";
			tmp(35,39) := "10001011";
			tmp(35,40) := "10000001";
			tmp(35,41) := "10000010";
			tmp(35,42) := "10000001";
			tmp(35,43) := "01110010";
			tmp(35,44) := "01100110";
			tmp(35,45) := "01101000";
			tmp(35,46) := "01101110";
			tmp(35,47) := "01101010";
			tmp(35,48) := "01100011";
			tmp(35,49) := "01101101";
			tmp(35,50) := "01101111";
			tmp(35,51) := "01110000";
			tmp(35,52) := "01100100";
			tmp(35,53) := "01011100";
			tmp(35,54) := "01011010";
			tmp(35,55) := "01010011";
			tmp(35,56) := "01001101";
			tmp(35,57) := "01010101";
			tmp(35,58) := "01010001";
			tmp(35,59) := "01010111";
			tmp(35,60) := "01101011";
			tmp(35,61) := "01111110";
			tmp(35,62) := "10001011";
			tmp(35,63) := "10000110";
			tmp(35,64) := "10000011";
			tmp(35,65) := "10001001";
			tmp(35,66) := "10001001";
			tmp(35,67) := "10001010";
			tmp(35,68) := "10000110";
			tmp(35,69) := "01110111";
			tmp(35,70) := "01111000";
			tmp(35,71) := "10001101";
			tmp(35,72) := "10010000";
			tmp(35,73) := "01111011";
			tmp(35,74) := "01110001";
			tmp(35,75) := "01111101";
			tmp(35,76) := "10000111";
			tmp(35,77) := "10000101";
			tmp(35,78) := "10110110";
			tmp(35,79) := "11110101";
			tmp(35,80) := "11111100";
			tmp(36,1) := "11111111";
			tmp(36,2) := "11111111";
			tmp(36,3) := "11111111";
			tmp(36,4) := "11111111";
			tmp(36,5) := "11111111";
			tmp(36,6) := "11111111";
			tmp(36,7) := "11111111";
			tmp(36,8) := "11111111";
			tmp(36,9) := "11111111";
			tmp(36,10) := "11111110";
			tmp(36,11) := "11111111";
			tmp(36,12) := "11111111";
			tmp(36,13) := "11111000";
			tmp(36,14) := "11101100";
			tmp(36,15) := "10101000";
			tmp(36,16) := "10110111";
			tmp(36,17) := "11111111";
			tmp(36,18) := "11101011";
			tmp(36,19) := "11101010";
			tmp(36,20) := "11101110";
			tmp(36,21) := "11101110";
			tmp(36,22) := "11101010";
			tmp(36,23) := "11011110";
			tmp(36,24) := "11100000";
			tmp(36,25) := "11101001";
			tmp(36,26) := "11010010";
			tmp(36,27) := "11010010";
			tmp(36,28) := "11011001";
			tmp(36,29) := "11010111";
			tmp(36,30) := "11000001";
			tmp(36,31) := "10111100";
			tmp(36,32) := "10111010";
			tmp(36,33) := "11001100";
			tmp(36,34) := "10110111";
			tmp(36,35) := "10101001";
			tmp(36,36) := "10010111";
			tmp(36,37) := "10001000";
			tmp(36,38) := "10001110";
			tmp(36,39) := "10000110";
			tmp(36,40) := "01111101";
			tmp(36,41) := "01111011";
			tmp(36,42) := "01111000";
			tmp(36,43) := "01101011";
			tmp(36,44) := "01101101";
			tmp(36,45) := "01110101";
			tmp(36,46) := "01110000";
			tmp(36,47) := "01100111";
			tmp(36,48) := "01101010";
			tmp(36,49) := "01110100";
			tmp(36,50) := "01110110";
			tmp(36,51) := "01101100";
			tmp(36,52) := "01101000";
			tmp(36,53) := "01100101";
			tmp(36,54) := "01011011";
			tmp(36,55) := "01010100";
			tmp(36,56) := "01001111";
			tmp(36,57) := "01010110";
			tmp(36,58) := "01100100";
			tmp(36,59) := "01101011";
			tmp(36,60) := "01110111";
			tmp(36,61) := "01111101";
			tmp(36,62) := "10000110";
			tmp(36,63) := "10001100";
			tmp(36,64) := "10001001";
			tmp(36,65) := "10010001";
			tmp(36,66) := "01111011";
			tmp(36,67) := "01111100";
			tmp(36,68) := "10000110";
			tmp(36,69) := "01111111";
			tmp(36,70) := "01111000";
			tmp(36,71) := "10000010";
			tmp(36,72) := "10000110";
			tmp(36,73) := "10000111";
			tmp(36,74) := "10000100";
			tmp(36,75) := "01111010";
			tmp(36,76) := "01111111";
			tmp(36,77) := "10001011";
			tmp(36,78) := "11010110";
			tmp(36,79) := "11110111";
			tmp(36,80) := "11111111";
			tmp(37,1) := "11111111";
			tmp(37,2) := "11111111";
			tmp(37,3) := "11111111";
			tmp(37,4) := "11111111";
			tmp(37,5) := "11111111";
			tmp(37,6) := "11111111";
			tmp(37,7) := "11111111";
			tmp(37,8) := "11111111";
			tmp(37,9) := "11111111";
			tmp(37,10) := "11111111";
			tmp(37,11) := "11111101";
			tmp(37,12) := "11111111";
			tmp(37,13) := "11111111";
			tmp(37,14) := "11111000";
			tmp(37,15) := "11001010";
			tmp(37,16) := "11110000";
			tmp(37,17) := "11110100";
			tmp(37,18) := "11110011";
			tmp(37,19) := "11101110";
			tmp(37,20) := "11011110";
			tmp(37,21) := "11100000";
			tmp(37,22) := "11011010";
			tmp(37,23) := "11001100";
			tmp(37,24) := "11001100";
			tmp(37,25) := "11010101";
			tmp(37,26) := "11010100";
			tmp(37,27) := "11011001";
			tmp(37,28) := "11100101";
			tmp(37,29) := "11100000";
			tmp(37,30) := "11001110";
			tmp(37,31) := "10111010";
			tmp(37,32) := "11000111";
			tmp(37,33) := "11010111";
			tmp(37,34) := "10110011";
			tmp(37,35) := "10101000";
			tmp(37,36) := "10011001";
			tmp(37,37) := "10010000";
			tmp(37,38) := "10001000";
			tmp(37,39) := "10000111";
			tmp(37,40) := "10000110";
			tmp(37,41) := "01111010";
			tmp(37,42) := "01110111";
			tmp(37,43) := "01101111";
			tmp(37,44) := "01110001";
			tmp(37,45) := "01110000";
			tmp(37,46) := "01101100";
			tmp(37,47) := "01110001";
			tmp(37,48) := "10000101";
			tmp(37,49) := "01110101";
			tmp(37,50) := "01110001";
			tmp(37,51) := "01101000";
			tmp(37,52) := "01100011";
			tmp(37,53) := "01011110";
			tmp(37,54) := "01010000";
			tmp(37,55) := "01001001";
			tmp(37,56) := "01000111";
			tmp(37,57) := "01100001";
			tmp(37,58) := "01110101";
			tmp(37,59) := "10000000";
			tmp(37,60) := "10000101";
			tmp(37,61) := "10000010";
			tmp(37,62) := "10001000";
			tmp(37,63) := "10010000";
			tmp(37,64) := "10010000";
			tmp(37,65) := "10001010";
			tmp(37,66) := "01111101";
			tmp(37,67) := "01110101";
			tmp(37,68) := "01110010";
			tmp(37,69) := "01111010";
			tmp(37,70) := "01111011";
			tmp(37,71) := "01110110";
			tmp(37,72) := "01111000";
			tmp(37,73) := "10000000";
			tmp(37,74) := "10001100";
			tmp(37,75) := "10001101";
			tmp(37,76) := "10001000";
			tmp(37,77) := "10100001";
			tmp(37,78) := "11011010";
			tmp(37,79) := "11111110";
			tmp(37,80) := "11111111";
			tmp(38,1) := "11111111";
			tmp(38,2) := "11111111";
			tmp(38,3) := "11111111";
			tmp(38,4) := "11111111";
			tmp(38,5) := "11111111";
			tmp(38,6) := "11111111";
			tmp(38,7) := "11111111";
			tmp(38,8) := "11111111";
			tmp(38,9) := "11111000";
			tmp(38,10) := "11111111";
			tmp(38,11) := "11111110";
			tmp(38,12) := "11111110";
			tmp(38,13) := "11111100";
			tmp(38,14) := "11111111";
			tmp(38,15) := "11110111";
			tmp(38,16) := "11110101";
			tmp(38,17) := "11111011";
			tmp(38,18) := "11110110";
			tmp(38,19) := "11111011";
			tmp(38,20) := "11111000";
			tmp(38,21) := "11011000";
			tmp(38,22) := "11010001";
			tmp(38,23) := "11010111";
			tmp(38,24) := "11011010";
			tmp(38,25) := "11011111";
			tmp(38,26) := "11011000";
			tmp(38,27) := "11001111";
			tmp(38,28) := "11100111";
			tmp(38,29) := "11100100";
			tmp(38,30) := "11000111";
			tmp(38,31) := "11000000";
			tmp(38,32) := "11000011";
			tmp(38,33) := "11001001";
			tmp(38,34) := "10101110";
			tmp(38,35) := "10100001";
			tmp(38,36) := "10010101";
			tmp(38,37) := "10010101";
			tmp(38,38) := "10001101";
			tmp(38,39) := "10010111";
			tmp(38,40) := "10000101";
			tmp(38,41) := "01111010";
			tmp(38,42) := "01110111";
			tmp(38,43) := "01110010";
			tmp(38,44) := "01110011";
			tmp(38,45) := "01101110";
			tmp(38,46) := "01110000";
			tmp(38,47) := "01110100";
			tmp(38,48) := "01111001";
			tmp(38,49) := "01111001";
			tmp(38,50) := "01101111";
			tmp(38,51) := "01101110";
			tmp(38,52) := "01100011";
			tmp(38,53) := "01010000";
			tmp(38,54) := "01001011";
			tmp(38,55) := "01001110";
			tmp(38,56) := "01011001";
			tmp(38,57) := "01011100";
			tmp(38,58) := "01110100";
			tmp(38,59) := "01111110";
			tmp(38,60) := "10001010";
			tmp(38,61) := "10000110";
			tmp(38,62) := "10001000";
			tmp(38,63) := "10001111";
			tmp(38,64) := "10001000";
			tmp(38,65) := "01111101";
			tmp(38,66) := "01111001";
			tmp(38,67) := "01101110";
			tmp(38,68) := "01101100";
			tmp(38,69) := "10000010";
			tmp(38,70) := "01111101";
			tmp(38,71) := "01101000";
			tmp(38,72) := "01110010";
			tmp(38,73) := "01110101";
			tmp(38,74) := "01111101";
			tmp(38,75) := "10001000";
			tmp(38,76) := "10001110";
			tmp(38,77) := "10101000";
			tmp(38,78) := "11111100";
			tmp(38,79) := "11111111";
			tmp(38,80) := "11111110";
			tmp(39,1) := "11111111";
			tmp(39,2) := "11111111";
			tmp(39,3) := "11111111";
			tmp(39,4) := "11111111";
			tmp(39,5) := "11111111";
			tmp(39,6) := "11111111";
			tmp(39,7) := "11111111";
			tmp(39,8) := "11111111";
			tmp(39,9) := "11111111";
			tmp(39,10) := "11111111";
			tmp(39,11) := "11111111";
			tmp(39,12) := "11111101";
			tmp(39,13) := "11111110";
			tmp(39,14) := "11111111";
			tmp(39,15) := "11111011";
			tmp(39,16) := "11111001";
			tmp(39,17) := "11100101";
			tmp(39,18) := "11100110";
			tmp(39,19) := "11100111";
			tmp(39,20) := "11011110";
			tmp(39,21) := "11010110";
			tmp(39,22) := "11010111";
			tmp(39,23) := "11001110";
			tmp(39,24) := "11010100";
			tmp(39,25) := "11101110";
			tmp(39,26) := "11100110";
			tmp(39,27) := "11001111";
			tmp(39,28) := "11011001";
			tmp(39,29) := "11001100";
			tmp(39,30) := "11000000";
			tmp(39,31) := "10110110";
			tmp(39,32) := "10111101";
			tmp(39,33) := "11000011";
			tmp(39,34) := "10101011";
			tmp(39,35) := "10100011";
			tmp(39,36) := "10110010";
			tmp(39,37) := "10100001";
			tmp(39,38) := "10011010";
			tmp(39,39) := "10011010";
			tmp(39,40) := "10001001";
			tmp(39,41) := "10000011";
			tmp(39,42) := "01111110";
			tmp(39,43) := "01110111";
			tmp(39,44) := "01110110";
			tmp(39,45) := "01110000";
			tmp(39,46) := "01110100";
			tmp(39,47) := "01110111";
			tmp(39,48) := "01110111";
			tmp(39,49) := "01111000";
			tmp(39,50) := "01101000";
			tmp(39,51) := "01100111";
			tmp(39,52) := "01100000";
			tmp(39,53) := "01010010";
			tmp(39,54) := "01001111";
			tmp(39,55) := "01010010";
			tmp(39,56) := "01100000";
			tmp(39,57) := "01101001";
			tmp(39,58) := "01110101";
			tmp(39,59) := "10000111";
			tmp(39,60) := "10001001";
			tmp(39,61) := "10000010";
			tmp(39,62) := "10000100";
			tmp(39,63) := "01111010";
			tmp(39,64) := "01111100";
			tmp(39,65) := "01111000";
			tmp(39,66) := "01101111";
			tmp(39,67) := "01101010";
			tmp(39,68) := "01101011";
			tmp(39,69) := "01111101";
			tmp(39,70) := "01111110";
			tmp(39,71) := "01110001";
			tmp(39,72) := "01101111";
			tmp(39,73) := "01101011";
			tmp(39,74) := "01101100";
			tmp(39,75) := "01111001";
			tmp(39,76) := "01111110";
			tmp(39,77) := "11000011";
			tmp(39,78) := "11111001";
			tmp(39,79) := "11111101";
			tmp(39,80) := "11111100";
			tmp(40,1) := "11111111";
			tmp(40,2) := "11111111";
			tmp(40,3) := "11111111";
			tmp(40,4) := "11111111";
			tmp(40,5) := "11111111";
			tmp(40,6) := "11111111";
			tmp(40,7) := "11111111";
			tmp(40,8) := "11111111";
			tmp(40,9) := "11111111";
			tmp(40,10) := "11111100";
			tmp(40,11) := "11111111";
			tmp(40,12) := "11111111";
			tmp(40,13) := "11111111";
			tmp(40,14) := "11111111";
			tmp(40,15) := "11111010";
			tmp(40,16) := "11101101";
			tmp(40,17) := "11101110";
			tmp(40,18) := "11011010";
			tmp(40,19) := "11011111";
			tmp(40,20) := "11011110";
			tmp(40,21) := "11011111";
			tmp(40,22) := "11100010";
			tmp(40,23) := "11011110";
			tmp(40,24) := "11100001";
			tmp(40,25) := "11100011";
			tmp(40,26) := "11011010";
			tmp(40,27) := "11100010";
			tmp(40,28) := "11011100";
			tmp(40,29) := "11010110";
			tmp(40,30) := "10111101";
			tmp(40,31) := "10111111";
			tmp(40,32) := "11001100";
			tmp(40,33) := "10111010";
			tmp(40,34) := "10100101";
			tmp(40,35) := "10100000";
			tmp(40,36) := "10010111";
			tmp(40,37) := "10100111";
			tmp(40,38) := "10010111";
			tmp(40,39) := "10001001";
			tmp(40,40) := "10000111";
			tmp(40,41) := "10000110";
			tmp(40,42) := "10000100";
			tmp(40,43) := "01111001";
			tmp(40,44) := "01110010";
			tmp(40,45) := "01111001";
			tmp(40,46) := "10000010";
			tmp(40,47) := "01111110";
			tmp(40,48) := "01110000";
			tmp(40,49) := "01101110";
			tmp(40,50) := "01100100";
			tmp(40,51) := "01100000";
			tmp(40,52) := "01011010";
			tmp(40,53) := "01001101";
			tmp(40,54) := "01001010";
			tmp(40,55) := "01100001";
			tmp(40,56) := "10000110";
			tmp(40,57) := "10000000";
			tmp(40,58) := "10000110";
			tmp(40,59) := "10000111";
			tmp(40,60) := "10001001";
			tmp(40,61) := "10000010";
			tmp(40,62) := "01111110";
			tmp(40,63) := "01110111";
			tmp(40,64) := "01101101";
			tmp(40,65) := "01110001";
			tmp(40,66) := "01111011";
			tmp(40,67) := "01110110";
			tmp(40,68) := "01101010";
			tmp(40,69) := "01101100";
			tmp(40,70) := "01101111";
			tmp(40,71) := "01110111";
			tmp(40,72) := "01111111";
			tmp(40,73) := "01110110";
			tmp(40,74) := "01101011";
			tmp(40,75) := "01111100";
			tmp(40,76) := "10100111";
			tmp(40,77) := "11111001";
			tmp(40,78) := "11111110";
			tmp(40,79) := "11111111";
			tmp(40,80) := "11111111";
			tmp(41,1) := "11111111";
			tmp(41,2) := "11111101";
			tmp(41,3) := "11111111";
			tmp(41,4) := "11111111";
			tmp(41,5) := "11111111";
			tmp(41,6) := "11111111";
			tmp(41,7) := "11111111";
			tmp(41,8) := "11111110";
			tmp(41,9) := "11111110";
			tmp(41,10) := "11111100";
			tmp(41,11) := "11111111";
			tmp(41,12) := "11111110";
			tmp(41,13) := "11111111";
			tmp(41,14) := "11111001";
			tmp(41,15) := "11111111";
			tmp(41,16) := "11110001";
			tmp(41,17) := "11011101";
			tmp(41,18) := "11100110";
			tmp(41,19) := "11100100";
			tmp(41,20) := "11011100";
			tmp(41,21) := "11100101";
			tmp(41,22) := "11011011";
			tmp(41,23) := "11010110";
			tmp(41,24) := "11001111";
			tmp(41,25) := "11011110";
			tmp(41,26) := "11101110";
			tmp(41,27) := "11101100";
			tmp(41,28) := "11101000";
			tmp(41,29) := "11010000";
			tmp(41,30) := "11000100";
			tmp(41,31) := "11000011";
			tmp(41,32) := "10111011";
			tmp(41,33) := "10101110";
			tmp(41,34) := "10110101";
			tmp(41,35) := "10100110";
			tmp(41,36) := "10011110";
			tmp(41,37) := "10010110";
			tmp(41,38) := "10010000";
			tmp(41,39) := "10011101";
			tmp(41,40) := "10001011";
			tmp(41,41) := "10000000";
			tmp(41,42) := "10001010";
			tmp(41,43) := "01111110";
			tmp(41,44) := "01110010";
			tmp(41,45) := "01111100";
			tmp(41,46) := "10010010";
			tmp(41,47) := "01111101";
			tmp(41,48) := "01101100";
			tmp(41,49) := "01100101";
			tmp(41,50) := "01011110";
			tmp(41,51) := "01010101";
			tmp(41,52) := "01001010";
			tmp(41,53) := "01001110";
			tmp(41,54) := "01010111";
			tmp(41,55) := "01100101";
			tmp(41,56) := "01111000";
			tmp(41,57) := "10001000";
			tmp(41,58) := "10000010";
			tmp(41,59) := "10000110";
			tmp(41,60) := "10001001";
			tmp(41,61) := "10000111";
			tmp(41,62) := "01111011";
			tmp(41,63) := "01111011";
			tmp(41,64) := "01110101";
			tmp(41,65) := "01110010";
			tmp(41,66) := "01101010";
			tmp(41,67) := "01101010";
			tmp(41,68) := "01100111";
			tmp(41,69) := "01100111";
			tmp(41,70) := "01100000";
			tmp(41,71) := "01110100";
			tmp(41,72) := "01111101";
			tmp(41,73) := "01111100";
			tmp(41,74) := "10000101";
			tmp(41,75) := "10000101";
			tmp(41,76) := "11001100";
			tmp(41,77) := "11111001";
			tmp(41,78) := "11111110";
			tmp(41,79) := "11111111";
			tmp(41,80) := "11111111";
			tmp(42,1) := "11111100";
			tmp(42,2) := "11111111";
			tmp(42,3) := "11111111";
			tmp(42,4) := "11111111";
			tmp(42,5) := "11111111";
			tmp(42,6) := "11111100";
			tmp(42,7) := "11111111";
			tmp(42,8) := "11111111";
			tmp(42,9) := "11111111";
			tmp(42,10) := "11111100";
			tmp(42,11) := "11111111";
			tmp(42,12) := "11111000";
			tmp(42,13) := "11111001";
			tmp(42,14) := "11111111";
			tmp(42,15) := "11111100";
			tmp(42,16) := "11110101";
			tmp(42,17) := "11011000";
			tmp(42,18) := "11100001";
			tmp(42,19) := "11010101";
			tmp(42,20) := "11011001";
			tmp(42,21) := "11010011";
			tmp(42,22) := "11010110";
			tmp(42,23) := "11010100";
			tmp(42,24) := "11000011";
			tmp(42,25) := "11001110";
			tmp(42,26) := "11011011";
			tmp(42,27) := "11010111";
			tmp(42,28) := "11001111";
			tmp(42,29) := "11001001";
			tmp(42,30) := "10111101";
			tmp(42,31) := "10111110";
			tmp(42,32) := "10110111";
			tmp(42,33) := "10110111";
			tmp(42,34) := "10101101";
			tmp(42,35) := "10100001";
			tmp(42,36) := "10100000";
			tmp(42,37) := "10011100";
			tmp(42,38) := "10110101";
			tmp(42,39) := "10011011";
			tmp(42,40) := "10010100";
			tmp(42,41) := "10001110";
			tmp(42,42) := "10000110";
			tmp(42,43) := "10000000";
			tmp(42,44) := "10000000";
			tmp(42,45) := "01111011";
			tmp(42,46) := "01111011";
			tmp(42,47) := "01110110";
			tmp(42,48) := "01101110";
			tmp(42,49) := "01101100";
			tmp(42,50) := "01101100";
			tmp(42,51) := "01011000";
			tmp(42,52) := "01001001";
			tmp(42,53) := "01010000";
			tmp(42,54) := "01010110";
			tmp(42,55) := "01101000";
			tmp(42,56) := "10000110";
			tmp(42,57) := "10000101";
			tmp(42,58) := "01111100";
			tmp(42,59) := "01111100";
			tmp(42,60) := "10000100";
			tmp(42,61) := "01111111";
			tmp(42,62) := "01111110";
			tmp(42,63) := "10000010";
			tmp(42,64) := "01110111";
			tmp(42,65) := "01101110";
			tmp(42,66) := "01100011";
			tmp(42,67) := "01100101";
			tmp(42,68) := "01110110";
			tmp(42,69) := "01100111";
			tmp(42,70) := "01101001";
			tmp(42,71) := "01100010";
			tmp(42,72) := "01011111";
			tmp(42,73) := "01110011";
			tmp(42,74) := "10000100";
			tmp(42,75) := "10011110";
			tmp(42,76) := "11110110";
			tmp(42,77) := "11111111";
			tmp(42,78) := "11111110";
			tmp(42,79) := "11111111";
			tmp(42,80) := "11111010";
			tmp(43,1) := "11111111";
			tmp(43,2) := "11111111";
			tmp(43,3) := "11111110";
			tmp(43,4) := "11111110";
			tmp(43,5) := "11111110";
			tmp(43,6) := "11111110";
			tmp(43,7) := "11111101";
			tmp(43,8) := "11110100";
			tmp(43,9) := "11011100";
			tmp(43,10) := "10111111";
			tmp(43,11) := "10010100";
			tmp(43,12) := "01100000";
			tmp(43,13) := "10000100";
			tmp(43,14) := "10101011";
			tmp(43,15) := "11100110";
			tmp(43,16) := "11101000";
			tmp(43,17) := "11011010";
			tmp(43,18) := "11000010";
			tmp(43,19) := "11001001";
			tmp(43,20) := "11000101";
			tmp(43,21) := "11001100";
			tmp(43,22) := "11011001";
			tmp(43,23) := "11100011";
			tmp(43,24) := "11011111";
			tmp(43,25) := "11001010";
			tmp(43,26) := "11010000";
			tmp(43,27) := "11010001";
			tmp(43,28) := "11011110";
			tmp(43,29) := "11001110";
			tmp(43,30) := "11000000";
			tmp(43,31) := "10111010";
			tmp(43,32) := "10110101";
			tmp(43,33) := "11000110";
			tmp(43,34) := "11010000";
			tmp(43,35) := "10110001";
			tmp(43,36) := "10100000";
			tmp(43,37) := "10100111";
			tmp(43,38) := "10110100";
			tmp(43,39) := "10100110";
			tmp(43,40) := "10010000";
			tmp(43,41) := "10010011";
			tmp(43,42) := "10001011";
			tmp(43,43) := "10000001";
			tmp(43,44) := "01111001";
			tmp(43,45) := "01111010";
			tmp(43,46) := "01110111";
			tmp(43,47) := "01110111";
			tmp(43,48) := "01101111";
			tmp(43,49) := "01101110";
			tmp(43,50) := "01011111";
			tmp(43,51) := "01010001";
			tmp(43,52) := "01010110";
			tmp(43,53) := "01100001";
			tmp(43,54) := "01100111";
			tmp(43,55) := "01110100";
			tmp(43,56) := "01111000";
			tmp(43,57) := "01110111";
			tmp(43,58) := "01111111";
			tmp(43,59) := "10000100";
			tmp(43,60) := "10001111";
			tmp(43,61) := "10000110";
			tmp(43,62) := "01111010";
			tmp(43,63) := "01101110";
			tmp(43,64) := "01110101";
			tmp(43,65) := "01101011";
			tmp(43,66) := "01101000";
			tmp(43,67) := "01101100";
			tmp(43,68) := "01111000";
			tmp(43,69) := "01110100";
			tmp(43,70) := "01110010";
			tmp(43,71) := "01101001";
			tmp(43,72) := "01110110";
			tmp(43,73) := "01101110";
			tmp(43,74) := "10000110";
			tmp(43,75) := "11001101";
			tmp(43,76) := "11111000";
			tmp(43,77) := "11111111";
			tmp(43,78) := "11111110";
			tmp(43,79) := "11111110";
			tmp(43,80) := "11111011";
			tmp(44,1) := "11111111";
			tmp(44,2) := "11111111";
			tmp(44,3) := "11111011";
			tmp(44,4) := "11111011";
			tmp(44,5) := "11111111";
			tmp(44,6) := "11111111";
			tmp(44,7) := "11011010";
			tmp(44,8) := "10100101";
			tmp(44,9) := "01100111";
			tmp(44,10) := "01000010";
			tmp(44,11) := "00111111";
			tmp(44,12) := "01001000";
			tmp(44,13) := "01010011";
			tmp(44,14) := "01001111";
			tmp(44,15) := "01010111";
			tmp(44,16) := "10000001";
			tmp(44,17) := "10101000";
			tmp(44,18) := "10110101";
			tmp(44,19) := "10110101";
			tmp(44,20) := "10110000";
			tmp(44,21) := "11000110";
			tmp(44,22) := "11100111";
			tmp(44,23) := "11101101";
			tmp(44,24) := "11011111";
			tmp(44,25) := "11100011";
			tmp(44,26) := "11100010";
			tmp(44,27) := "11010100";
			tmp(44,28) := "11011001";
			tmp(44,29) := "11011010";
			tmp(44,30) := "11000110";
			tmp(44,31) := "10111100";
			tmp(44,32) := "11000000";
			tmp(44,33) := "11011011";
			tmp(44,34) := "11010101";
			tmp(44,35) := "10110011";
			tmp(44,36) := "10100101";
			tmp(44,37) := "10101010";
			tmp(44,38) := "10100011";
			tmp(44,39) := "10011000";
			tmp(44,40) := "10010001";
			tmp(44,41) := "10001011";
			tmp(44,42) := "10000101";
			tmp(44,43) := "01111100";
			tmp(44,44) := "01110100";
			tmp(44,45) := "01110011";
			tmp(44,46) := "01101110";
			tmp(44,47) := "01101010";
			tmp(44,48) := "01100111";
			tmp(44,49) := "01011000";
			tmp(44,50) := "01001011";
			tmp(44,51) := "01010101";
			tmp(44,52) := "01011011";
			tmp(44,53) := "01110001";
			tmp(44,54) := "10000001";
			tmp(44,55) := "01111100";
			tmp(44,56) := "10001001";
			tmp(44,57) := "01111111";
			tmp(44,58) := "01111000";
			tmp(44,59) := "01111101";
			tmp(44,60) := "10001011";
			tmp(44,61) := "10001001";
			tmp(44,62) := "01111000";
			tmp(44,63) := "01100100";
			tmp(44,64) := "01101110";
			tmp(44,65) := "01110011";
			tmp(44,66) := "01111000";
			tmp(44,67) := "01100010";
			tmp(44,68) := "01100010";
			tmp(44,69) := "01100111";
			tmp(44,70) := "01100111";
			tmp(44,71) := "01110111";
			tmp(44,72) := "10000001";
			tmp(44,73) := "10010101";
			tmp(44,74) := "11001111";
			tmp(44,75) := "11111111";
			tmp(44,76) := "11111100";
			tmp(44,77) := "11111110";
			tmp(44,78) := "11111111";
			tmp(44,79) := "11111110";
			tmp(44,80) := "11111111";
			tmp(45,1) := "11111111";
			tmp(45,2) := "11111111";
			tmp(45,3) := "11111011";
			tmp(45,4) := "11111111";
			tmp(45,5) := "11110101";
			tmp(45,6) := "11001011";
			tmp(45,7) := "10000000";
			tmp(45,8) := "01001010";
			tmp(45,9) := "00110111";
			tmp(45,10) := "01000000";
			tmp(45,11) := "01001100";
			tmp(45,12) := "01000101";
			tmp(45,13) := "01001011";
			tmp(45,14) := "01001010";
			tmp(45,15) := "01001001";
			tmp(45,16) := "01000110";
			tmp(45,17) := "01101001";
			tmp(45,18) := "10100001";
			tmp(45,19) := "10011101";
			tmp(45,20) := "10100100";
			tmp(45,21) := "10111100";
			tmp(45,22) := "11001110";
			tmp(45,23) := "11011111";
			tmp(45,24) := "11011100";
			tmp(45,25) := "11011011";
			tmp(45,26) := "11010001";
			tmp(45,27) := "11010100";
			tmp(45,28) := "11100001";
			tmp(45,29) := "11101011";
			tmp(45,30) := "11011001";
			tmp(45,31) := "10111110";
			tmp(45,32) := "10110111";
			tmp(45,33) := "11000100";
			tmp(45,34) := "11001001";
			tmp(45,35) := "10110111";
			tmp(45,36) := "10100110";
			tmp(45,37) := "10011010";
			tmp(45,38) := "10001011";
			tmp(45,39) := "10011100";
			tmp(45,40) := "10001110";
			tmp(45,41) := "10001011";
			tmp(45,42) := "01111110";
			tmp(45,43) := "01111010";
			tmp(45,44) := "10000010";
			tmp(45,45) := "01111011";
			tmp(45,46) := "01111010";
			tmp(45,47) := "01110011";
			tmp(45,48) := "01011011";
			tmp(45,49) := "01001111";
			tmp(45,50) := "01011000";
			tmp(45,51) := "01101000";
			tmp(45,52) := "01110001";
			tmp(45,53) := "10000100";
			tmp(45,54) := "10010010";
			tmp(45,55) := "01111111";
			tmp(45,56) := "01110111";
			tmp(45,57) := "01111010";
			tmp(45,58) := "01111001";
			tmp(45,59) := "01111101";
			tmp(45,60) := "01111110";
			tmp(45,61) := "10000001";
			tmp(45,62) := "01111101";
			tmp(45,63) := "01110011";
			tmp(45,64) := "01101110";
			tmp(45,65) := "01101111";
			tmp(45,66) := "01111101";
			tmp(45,67) := "01100011";
			tmp(45,68) := "01101100";
			tmp(45,69) := "01100111";
			tmp(45,70) := "01101001";
			tmp(45,71) := "01111001";
			tmp(45,72) := "10001101";
			tmp(45,73) := "10110101";
			tmp(45,74) := "11101010";
			tmp(45,75) := "11111010";
			tmp(45,76) := "11111110";
			tmp(45,77) := "11111010";
			tmp(45,78) := "11111101";
			tmp(45,79) := "11111110";
			tmp(45,80) := "11111111";
			tmp(46,1) := "11111110";
			tmp(46,2) := "11111111";
			tmp(46,3) := "11111111";
			tmp(46,4) := "11111101";
			tmp(46,5) := "11000101";
			tmp(46,6) := "01100101";
			tmp(46,7) := "00110101";
			tmp(46,8) := "00110101";
			tmp(46,9) := "01000000";
			tmp(46,10) := "01000111";
			tmp(46,11) := "01001010";
			tmp(46,12) := "01000111";
			tmp(46,13) := "01000101";
			tmp(46,14) := "01001101";
			tmp(46,15) := "01001011";
			tmp(46,16) := "01001010";
			tmp(46,17) := "01011000";
			tmp(46,18) := "01111100";
			tmp(46,19) := "10010101";
			tmp(46,20) := "10001101";
			tmp(46,21) := "10011101";
			tmp(46,22) := "11000011";
			tmp(46,23) := "11100011";
			tmp(46,24) := "11110010";
			tmp(46,25) := "11100101";
			tmp(46,26) := "11010100";
			tmp(46,27) := "11010101";
			tmp(46,28) := "11001010";
			tmp(46,29) := "11001101";
			tmp(46,30) := "11000100";
			tmp(46,31) := "11001010";
			tmp(46,32) := "11000000";
			tmp(46,33) := "10111000";
			tmp(46,34) := "10110101";
			tmp(46,35) := "10110101";
			tmp(46,36) := "10100100";
			tmp(46,37) := "10110000";
			tmp(46,38) := "10100010";
			tmp(46,39) := "10010011";
			tmp(46,40) := "10001101";
			tmp(46,41) := "10000101";
			tmp(46,42) := "10001100";
			tmp(46,43) := "01110101";
			tmp(46,44) := "01101101";
			tmp(46,45) := "01101111";
			tmp(46,46) := "01101101";
			tmp(46,47) := "01100101";
			tmp(46,48) := "01011100";
			tmp(46,49) := "01011001";
			tmp(46,50) := "01100101";
			tmp(46,51) := "01101111";
			tmp(46,52) := "01111001";
			tmp(46,53) := "10001110";
			tmp(46,54) := "10001101";
			tmp(46,55) := "01101110";
			tmp(46,56) := "01110100";
			tmp(46,57) := "01110100";
			tmp(46,58) := "01110010";
			tmp(46,59) := "01110010";
			tmp(46,60) := "01111000";
			tmp(46,61) := "01111111";
			tmp(46,62) := "01111100";
			tmp(46,63) := "01110010";
			tmp(46,64) := "01011111";
			tmp(46,65) := "01110100";
			tmp(46,66) := "01110011";
			tmp(46,67) := "01110110";
			tmp(46,68) := "10000001";
			tmp(46,69) := "01111010";
			tmp(46,70) := "10000010";
			tmp(46,71) := "10000101";
			tmp(46,72) := "10111101";
			tmp(46,73) := "11110110";
			tmp(46,74) := "11111111";
			tmp(46,75) := "11111111";
			tmp(46,76) := "11111110";
			tmp(46,77) := "11111110";
			tmp(46,78) := "11111111";
			tmp(46,79) := "11111101";
			tmp(46,80) := "11111111";
			tmp(47,1) := "11111010";
			tmp(47,2) := "11111111";
			tmp(47,3) := "11111110";
			tmp(47,4) := "11000110";
			tmp(47,5) := "01000100";
			tmp(47,6) := "00101000";
			tmp(47,7) := "00110110";
			tmp(47,8) := "00111111";
			tmp(47,9) := "00111101";
			tmp(47,10) := "00111111";
			tmp(47,11) := "01000011";
			tmp(47,12) := "01001010";
			tmp(47,13) := "01001101";
			tmp(47,14) := "01001110";
			tmp(47,15) := "01001000";
			tmp(47,16) := "01001010";
			tmp(47,17) := "01010101";
			tmp(47,18) := "01101010";
			tmp(47,19) := "10001001";
			tmp(47,20) := "10010011";
			tmp(47,21) := "10000111";
			tmp(47,22) := "10100111";
			tmp(47,23) := "11001111";
			tmp(47,24) := "11100000";
			tmp(47,25) := "11100001";
			tmp(47,26) := "11010001";
			tmp(47,27) := "11000101";
			tmp(47,28) := "11010100";
			tmp(47,29) := "11001111";
			tmp(47,30) := "10111101";
			tmp(47,31) := "11000111";
			tmp(47,32) := "11001001";
			tmp(47,33) := "11101001";
			tmp(47,34) := "11000110";
			tmp(47,35) := "10110010";
			tmp(47,36) := "10101011";
			tmp(47,37) := "10100001";
			tmp(47,38) := "10100001";
			tmp(47,39) := "10011100";
			tmp(47,40) := "10001100";
			tmp(47,41) := "10001000";
			tmp(47,42) := "10000010";
			tmp(47,43) := "01110010";
			tmp(47,44) := "01101000";
			tmp(47,45) := "01100101";
			tmp(47,46) := "01100001";
			tmp(47,47) := "01011101";
			tmp(47,48) := "01011011";
			tmp(47,49) := "01101110";
			tmp(47,50) := "10000001";
			tmp(47,51) := "10000110";
			tmp(47,52) := "10000110";
			tmp(47,53) := "01111111";
			tmp(47,54) := "01111100";
			tmp(47,55) := "01111011";
			tmp(47,56) := "01110111";
			tmp(47,57) := "01110011";
			tmp(47,58) := "01101111";
			tmp(47,59) := "01110001";
			tmp(47,60) := "01101011";
			tmp(47,61) := "01100011";
			tmp(47,62) := "01110110";
			tmp(47,63) := "01111011";
			tmp(47,64) := "01101000";
			tmp(47,65) := "01101101";
			tmp(47,66) := "01101110";
			tmp(47,67) := "01110001";
			tmp(47,68) := "01111001";
			tmp(47,69) := "10000110";
			tmp(47,70) := "10010111";
			tmp(47,71) := "10111001";
			tmp(47,72) := "11110000";
			tmp(47,73) := "11111101";
			tmp(47,74) := "11111111";
			tmp(47,75) := "11111111";
			tmp(47,76) := "11111111";
			tmp(47,77) := "11111111";
			tmp(47,78) := "11111110";
			tmp(47,79) := "11111111";
			tmp(47,80) := "11111101";
			tmp(48,1) := "11111111";
			tmp(48,2) := "11110111";
			tmp(48,3) := "11010000";
			tmp(48,4) := "01011011";
			tmp(48,5) := "00110100";
			tmp(48,6) := "00110100";
			tmp(48,7) := "00111101";
			tmp(48,8) := "01000000";
			tmp(48,9) := "00111111";
			tmp(48,10) := "01000011";
			tmp(48,11) := "01000110";
			tmp(48,12) := "01000111";
			tmp(48,13) := "01000100";
			tmp(48,14) := "00101110";
			tmp(48,15) := "00101101";
			tmp(48,16) := "00110100";
			tmp(48,17) := "00101111";
			tmp(48,18) := "00111100";
			tmp(48,19) := "01100000";
			tmp(48,20) := "10001000";
			tmp(48,21) := "10000011";
			tmp(48,22) := "10000111";
			tmp(48,23) := "10101101";
			tmp(48,24) := "11001001";
			tmp(48,25) := "11010101";
			tmp(48,26) := "11001011";
			tmp(48,27) := "11001111";
			tmp(48,28) := "11011000";
			tmp(48,29) := "11001100";
			tmp(48,30) := "11001010";
			tmp(48,31) := "11000111";
			tmp(48,32) := "11000011";
			tmp(48,33) := "11000011";
			tmp(48,34) := "10110001";
			tmp(48,35) := "10110001";
			tmp(48,36) := "10100101";
			tmp(48,37) := "10011110";
			tmp(48,38) := "10010011";
			tmp(48,39) := "10010110";
			tmp(48,40) := "01111101";
			tmp(48,41) := "01101100";
			tmp(48,42) := "01101010";
			tmp(48,43) := "01101100";
			tmp(48,44) := "01011011";
			tmp(48,45) := "01100111";
			tmp(48,46) := "01101001";
			tmp(48,47) := "01101001";
			tmp(48,48) := "01111001";
			tmp(48,49) := "10011000";
			tmp(48,50) := "10010101";
			tmp(48,51) := "10010000";
			tmp(48,52) := "10001110";
			tmp(48,53) := "10000110";
			tmp(48,54) := "01111100";
			tmp(48,55) := "01110110";
			tmp(48,56) := "01111011";
			tmp(48,57) := "01110010";
			tmp(48,58) := "01101100";
			tmp(48,59) := "01110110";
			tmp(48,60) := "01111010";
			tmp(48,61) := "01101100";
			tmp(48,62) := "01110001";
			tmp(48,63) := "01101001";
			tmp(48,64) := "01110110";
			tmp(48,65) := "01101101";
			tmp(48,66) := "01100111";
			tmp(48,67) := "01110000";
			tmp(48,68) := "01111001";
			tmp(48,69) := "10011110";
			tmp(48,70) := "11001110";
			tmp(48,71) := "11110000";
			tmp(48,72) := "11111110";
			tmp(48,73) := "11111110";
			tmp(48,74) := "11111110";
			tmp(48,75) := "11111101";
			tmp(48,76) := "11111111";
			tmp(48,77) := "11111111";
			tmp(48,78) := "11111000";
			tmp(48,79) := "11111110";
			tmp(48,80) := "11111111";
			tmp(49,1) := "11111110";
			tmp(49,2) := "11101101";
			tmp(49,3) := "10000001";
			tmp(49,4) := "00110001";
			tmp(49,5) := "00111000";
			tmp(49,6) := "00110111";
			tmp(49,7) := "00110100";
			tmp(49,8) := "00110011";
			tmp(49,9) := "00110110";
			tmp(49,10) := "01000101";
			tmp(49,11) := "01010101";
			tmp(49,12) := "01011010";
			tmp(49,13) := "01010000";
			tmp(49,14) := "01000100";
			tmp(49,15) := "00111111";
			tmp(49,16) := "00111111";
			tmp(49,17) := "00111011";
			tmp(49,18) := "00111000";
			tmp(49,19) := "01000000";
			tmp(49,20) := "01010111";
			tmp(49,21) := "01101001";
			tmp(49,22) := "01101101";
			tmp(49,23) := "10001110";
			tmp(49,24) := "10110011";
			tmp(49,25) := "11000101";
			tmp(49,26) := "11001011";
			tmp(49,27) := "11010110";
			tmp(49,28) := "11001001";
			tmp(49,29) := "11000010";
			tmp(49,30) := "11001010";
			tmp(49,31) := "11000101";
			tmp(49,32) := "10110011";
			tmp(49,33) := "10111110";
			tmp(49,34) := "10101011";
			tmp(49,35) := "10100110";
			tmp(49,36) := "10100100";
			tmp(49,37) := "10010100";
			tmp(49,38) := "10010100";
			tmp(49,39) := "10001001";
			tmp(49,40) := "01111011";
			tmp(49,41) := "01110001";
			tmp(49,42) := "01110110";
			tmp(49,43) := "01101011";
			tmp(49,44) := "01101100";
			tmp(49,45) := "01110001";
			tmp(49,46) := "01111010";
			tmp(49,47) := "10000100";
			tmp(49,48) := "10000101";
			tmp(49,49) := "10001111";
			tmp(49,50) := "10010101";
			tmp(49,51) := "10001010";
			tmp(49,52) := "10001100";
			tmp(49,53) := "10001001";
			tmp(49,54) := "01111011";
			tmp(49,55) := "01100110";
			tmp(49,56) := "01110000";
			tmp(49,57) := "01110010";
			tmp(49,58) := "01110010";
			tmp(49,59) := "01111011";
			tmp(49,60) := "01110110";
			tmp(49,61) := "01111010";
			tmp(49,62) := "01110011";
			tmp(49,63) := "01100000";
			tmp(49,64) := "01110110";
			tmp(49,65) := "01110011";
			tmp(49,66) := "10010001";
			tmp(49,67) := "10000000";
			tmp(49,68) := "10011110";
			tmp(49,69) := "11011011";
			tmp(49,70) := "11111100";
			tmp(49,71) := "11111111";
			tmp(49,72) := "11111111";
			tmp(49,73) := "11111111";
			tmp(49,74) := "11111111";
			tmp(49,75) := "11111111";
			tmp(49,76) := "11111111";
			tmp(49,77) := "11111111";
			tmp(49,78) := "11111111";
			tmp(49,79) := "11111111";
			tmp(49,80) := "11111111";
			tmp(50,1) := "11110100";
			tmp(50,2) := "10010111";
			tmp(50,3) := "01000101";
			tmp(50,4) := "00110111";
			tmp(50,5) := "00110111";
			tmp(50,6) := "00111110";
			tmp(50,7) := "00111001";
			tmp(50,8) := "00111100";
			tmp(50,9) := "00111101";
			tmp(50,10) := "01010111";
			tmp(50,11) := "01010100";
			tmp(50,12) := "01001010";
			tmp(50,13) := "01001100";
			tmp(50,14) := "01001101";
			tmp(50,15) := "01000111";
			tmp(50,16) := "01001010";
			tmp(50,17) := "01000111";
			tmp(50,18) := "01000110";
			tmp(50,19) := "00111001";
			tmp(50,20) := "00110111";
			tmp(50,21) := "01000001";
			tmp(50,22) := "01010110";
			tmp(50,23) := "01110001";
			tmp(50,24) := "10010101";
			tmp(50,25) := "10101011";
			tmp(50,26) := "10111011";
			tmp(50,27) := "10111110";
			tmp(50,28) := "10110100";
			tmp(50,29) := "11001101";
			tmp(50,30) := "10110111";
			tmp(50,31) := "10111110";
			tmp(50,32) := "10111001";
			tmp(50,33) := "10100110";
			tmp(50,34) := "10111000";
			tmp(50,35) := "10011101";
			tmp(50,36) := "10010001";
			tmp(50,37) := "10011000";
			tmp(50,38) := "10001011";
			tmp(50,39) := "01111101";
			tmp(50,40) := "01110100";
			tmp(50,41) := "01101100";
			tmp(50,42) := "01110000";
			tmp(50,43) := "01101110";
			tmp(50,44) := "10000101";
			tmp(50,45) := "10010100";
			tmp(50,46) := "10000110";
			tmp(50,47) := "01111111";
			tmp(50,48) := "10001001";
			tmp(50,49) := "10001100";
			tmp(50,50) := "10010010";
			tmp(50,51) := "10100110";
			tmp(50,52) := "10011011";
			tmp(50,53) := "01111111";
			tmp(50,54) := "01110001";
			tmp(50,55) := "01101100";
			tmp(50,56) := "01100110";
			tmp(50,57) := "01100111";
			tmp(50,58) := "01100111";
			tmp(50,59) := "01101000";
			tmp(50,60) := "01110111";
			tmp(50,61) := "10011010";
			tmp(50,62) := "01110010";
			tmp(50,63) := "01101101";
			tmp(50,64) := "01110011";
			tmp(50,65) := "10001000";
			tmp(50,66) := "10100110";
			tmp(50,67) := "11010001";
			tmp(50,68) := "11100101";
			tmp(50,69) := "11111010";
			tmp(50,70) := "11111001";
			tmp(50,71) := "11111110";
			tmp(50,72) := "11111011";
			tmp(50,73) := "11111111";
			tmp(50,74) := "11111111";
			tmp(50,75) := "11111111";
			tmp(50,76) := "11111111";
			tmp(50,77) := "11111111";
			tmp(50,78) := "11111111";
			tmp(50,79) := "11111111";
			tmp(50,80) := "11111111";
			tmp(51,1) := "11100110";
			tmp(51,2) := "01110111";
			tmp(51,3) := "00110110";
			tmp(51,4) := "00101111";
			tmp(51,5) := "00110100";
			tmp(51,6) := "00111000";
			tmp(51,7) := "00110101";
			tmp(51,8) := "00110011";
			tmp(51,9) := "01010101";
			tmp(51,10) := "01100101";
			tmp(51,11) := "01001101";
			tmp(51,12) := "01001111";
			tmp(51,13) := "01001000";
			tmp(51,14) := "00111101";
			tmp(51,15) := "00111110";
			tmp(51,16) := "01000000";
			tmp(51,17) := "00111101";
			tmp(51,18) := "00110100";
			tmp(51,19) := "00101100";
			tmp(51,20) := "00110111";
			tmp(51,21) := "01000001";
			tmp(51,22) := "01000110";
			tmp(51,23) := "01011010";
			tmp(51,24) := "01111101";
			tmp(51,25) := "10000010";
			tmp(51,26) := "10011111";
			tmp(51,27) := "10110000";
			tmp(51,28) := "10111100";
			tmp(51,29) := "11001001";
			tmp(51,30) := "10111010";
			tmp(51,31) := "10110111";
			tmp(51,32) := "10110101";
			tmp(51,33) := "10110001";
			tmp(51,34) := "10101001";
			tmp(51,35) := "10100000";
			tmp(51,36) := "10001100";
			tmp(51,37) := "10000010";
			tmp(51,38) := "10000101";
			tmp(51,39) := "10000000";
			tmp(51,40) := "01111000";
			tmp(51,41) := "01110110";
			tmp(51,42) := "01110100";
			tmp(51,43) := "10000001";
			tmp(51,44) := "10011100";
			tmp(51,45) := "10100101";
			tmp(51,46) := "10100001";
			tmp(51,47) := "10010111";
			tmp(51,48) := "10001011";
			tmp(51,49) := "10000111";
			tmp(51,50) := "01111111";
			tmp(51,51) := "10011011";
			tmp(51,52) := "10011001";
			tmp(51,53) := "10001110";
			tmp(51,54) := "01110110";
			tmp(51,55) := "01110000";
			tmp(51,56) := "01101000";
			tmp(51,57) := "01100111";
			tmp(51,58) := "01111001";
			tmp(51,59) := "01101101";
			tmp(51,60) := "01110001";
			tmp(51,61) := "01111110";
			tmp(51,62) := "01110111";
			tmp(51,63) := "01101001";
			tmp(51,64) := "01111111";
			tmp(51,65) := "10010000";
			tmp(51,66) := "11100010";
			tmp(51,67) := "11111011";
			tmp(51,68) := "11111111";
			tmp(51,69) := "11111110";
			tmp(51,70) := "11111111";
			tmp(51,71) := "11111111";
			tmp(51,72) := "11111111";
			tmp(51,73) := "11111110";
			tmp(51,74) := "11111111";
			tmp(51,75) := "11111111";
			tmp(51,76) := "11111111";
			tmp(51,77) := "11111111";
			tmp(51,78) := "11111111";
			tmp(51,79) := "11111111";
			tmp(51,80) := "11111111";
			tmp(52,1) := "11111100";
			tmp(52,2) := "11010111";
			tmp(52,3) := "10011100";
			tmp(52,4) := "10000110";
			tmp(52,5) := "01111101";
			tmp(52,6) := "01010110";
			tmp(52,7) := "00110000";
			tmp(52,8) := "01000110";
			tmp(52,9) := "01110001";
			tmp(52,10) := "01010100";
			tmp(52,11) := "01000100";
			tmp(52,12) := "01000110";
			tmp(52,13) := "01010011";
			tmp(52,14) := "01011001";
			tmp(52,15) := "01010111";
			tmp(52,16) := "01100010";
			tmp(52,17) := "01100111";
			tmp(52,18) := "10010011";
			tmp(52,19) := "10111011";
			tmp(52,20) := "11010001";
			tmp(52,21) := "11100111";
			tmp(52,22) := "11011011";
			tmp(52,23) := "11011001";
			tmp(52,24) := "10010100";
			tmp(52,25) := "01110010";
			tmp(52,26) := "10010000";
			tmp(52,27) := "10110000";
			tmp(52,28) := "10101111";
			tmp(52,29) := "10111101";
			tmp(52,30) := "10101100";
			tmp(52,31) := "10101110";
			tmp(52,32) := "10101000";
			tmp(52,33) := "10011101";
			tmp(52,34) := "10011010";
			tmp(52,35) := "10010010";
			tmp(52,36) := "10001101";
			tmp(52,37) := "10001011";
			tmp(52,38) := "10000000";
			tmp(52,39) := "01110111";
			tmp(52,40) := "01111111";
			tmp(52,41) := "10001100";
			tmp(52,42) := "10010101";
			tmp(52,43) := "10010111";
			tmp(52,44) := "10010010";
			tmp(52,45) := "10011101";
			tmp(52,46) := "10100011";
			tmp(52,47) := "10011011";
			tmp(52,48) := "10011010";
			tmp(52,49) := "10001000";
			tmp(52,50) := "01111110";
			tmp(52,51) := "10001011";
			tmp(52,52) := "10001011";
			tmp(52,53) := "10000010";
			tmp(52,54) := "10000001";
			tmp(52,55) := "10000101";
			tmp(52,56) := "01110100";
			tmp(52,57) := "10000011";
			tmp(52,58) := "10000001";
			tmp(52,59) := "01110100";
			tmp(52,60) := "01111010";
			tmp(52,61) := "01101000";
			tmp(52,62) := "01111010";
			tmp(52,63) := "10000101";
			tmp(52,64) := "10111100";
			tmp(52,65) := "11110001";
			tmp(52,66) := "11111111";
			tmp(52,67) := "11111110";
			tmp(52,68) := "11111111";
			tmp(52,69) := "11111111";
			tmp(52,70) := "11111101";
			tmp(52,71) := "11111111";
			tmp(52,72) := "11111110";
			tmp(52,73) := "11111110";
			tmp(52,74) := "11111110";
			tmp(52,75) := "11111111";
			tmp(52,76) := "11111111";
			tmp(52,77) := "11111111";
			tmp(52,78) := "11111111";
			tmp(52,79) := "11111111";
			tmp(52,80) := "11111111";
			tmp(53,1) := "11111111";
			tmp(53,2) := "11111101";
			tmp(53,3) := "11111110";
			tmp(53,4) := "11111100";
			tmp(53,5) := "11011001";
			tmp(53,6) := "01101001";
			tmp(53,7) := "00111111";
			tmp(53,8) := "01101111";
			tmp(53,9) := "01110101";
			tmp(53,10) := "01010011";
			tmp(53,11) := "01000100";
			tmp(53,12) := "01001011";
			tmp(53,13) := "01001101";
			tmp(53,14) := "01010000";
			tmp(53,15) := "01011100";
			tmp(53,16) := "10001001";
			tmp(53,17) := "11010011";
			tmp(53,18) := "11111011";
			tmp(53,19) := "11111111";
			tmp(53,20) := "11111111";
			tmp(53,21) := "11111101";
			tmp(53,22) := "11111100";
			tmp(53,23) := "11111001";
			tmp(53,24) := "11010000";
			tmp(53,25) := "01110010";
			tmp(53,26) := "10001111";
			tmp(53,27) := "10011000";
			tmp(53,28) := "10100000";
			tmp(53,29) := "10011101";
			tmp(53,30) := "10011010";
			tmp(53,31) := "10011101";
			tmp(53,32) := "10011101";
			tmp(53,33) := "10001110";
			tmp(53,34) := "10001010";
			tmp(53,35) := "10000110";
			tmp(53,36) := "10000011";
			tmp(53,37) := "10001101";
			tmp(53,38) := "10010011";
			tmp(53,39) := "10101100";
			tmp(53,40) := "10110000";
			tmp(53,41) := "10010110";
			tmp(53,42) := "10100000";
			tmp(53,43) := "10101011";
			tmp(53,44) := "10011111";
			tmp(53,45) := "10011100";
			tmp(53,46) := "10100100";
			tmp(53,47) := "10011101";
			tmp(53,48) := "10011100";
			tmp(53,49) := "10000011";
			tmp(53,50) := "01110110";
			tmp(53,51) := "01110110";
			tmp(53,52) := "10000001";
			tmp(53,53) := "10000010";
			tmp(53,54) := "01110101";
			tmp(53,55) := "01111000";
			tmp(53,56) := "10000100";
			tmp(53,57) := "10001110";
			tmp(53,58) := "10000110";
			tmp(53,59) := "10101010";
			tmp(53,60) := "10000101";
			tmp(53,61) := "01111101";
			tmp(53,62) := "10010000";
			tmp(53,63) := "10111000";
			tmp(53,64) := "11110011";
			tmp(53,65) := "11111111";
			tmp(53,66) := "11111000";
			tmp(53,67) := "11111001";
			tmp(53,68) := "11111000";
			tmp(53,69) := "11111110";
			tmp(53,70) := "11111110";
			tmp(53,71) := "11111101";
			tmp(53,72) := "11111110";
			tmp(53,73) := "11111110";
			tmp(53,74) := "11111110";
			tmp(53,75) := "11111111";
			tmp(53,76) := "11111111";
			tmp(53,77) := "11111111";
			tmp(53,78) := "11111111";
			tmp(53,79) := "11111111";
			tmp(53,80) := "11111111";
			tmp(54,1) := "11111111";
			tmp(54,2) := "11111100";
			tmp(54,3) := "11111100";
			tmp(54,4) := "11101111";
			tmp(54,5) := "10000101";
			tmp(54,6) := "00101000";
			tmp(54,7) := "01001101";
			tmp(54,8) := "01111010";
			tmp(54,9) := "01011000";
			tmp(54,10) := "00111110";
			tmp(54,11) := "00110010";
			tmp(54,12) := "00110101";
			tmp(54,13) := "01001001";
			tmp(54,14) := "01101100";
			tmp(54,15) := "10101010";
			tmp(54,16) := "11100101";
			tmp(54,17) := "11111111";
			tmp(54,18) := "11111001";
			tmp(54,19) := "11111111";
			tmp(54,20) := "11111111";
			tmp(54,21) := "11111111";
			tmp(54,22) := "11111111";
			tmp(54,23) := "11110110";
			tmp(54,24) := "10100000";
			tmp(54,25) := "01100110";
			tmp(54,26) := "10010000";
			tmp(54,27) := "10011110";
			tmp(54,28) := "01101010";
			tmp(54,29) := "10001000";
			tmp(54,30) := "01111001";
			tmp(54,31) := "01111100";
			tmp(54,32) := "01111111";
			tmp(54,33) := "10000101";
			tmp(54,34) := "10100001";
			tmp(54,35) := "10101010";
			tmp(54,36) := "01111010";
			tmp(54,37) := "10001011";
			tmp(54,38) := "10100100";
			tmp(54,39) := "11000111";
			tmp(54,40) := "11010001";
			tmp(54,41) := "10100101";
			tmp(54,42) := "10100011";
			tmp(54,43) := "10100100";
			tmp(54,44) := "10011011";
			tmp(54,45) := "10100100";
			tmp(54,46) := "10110001";
			tmp(54,47) := "10100110";
			tmp(54,48) := "10011110";
			tmp(54,49) := "10001001";
			tmp(54,50) := "10000001";
			tmp(54,51) := "01111010";
			tmp(54,52) := "01110110";
			tmp(54,53) := "01110100";
			tmp(54,54) := "01111101";
			tmp(54,55) := "01101101";
			tmp(54,56) := "01111000";
			tmp(54,57) := "10001101";
			tmp(54,58) := "10011100";
			tmp(54,59) := "10010001";
			tmp(54,60) := "01110010";
			tmp(54,61) := "10100010";
			tmp(54,62) := "11010010";
			tmp(54,63) := "11100100";
			tmp(54,64) := "11111000";
			tmp(54,65) := "11111111";
			tmp(54,66) := "11111111";
			tmp(54,67) := "11111100";
			tmp(54,68) := "11111111";
			tmp(54,69) := "11111100";
			tmp(54,70) := "11111111";
			tmp(54,71) := "11111111";
			tmp(54,72) := "11111101";
			tmp(54,73) := "11111110";
			tmp(54,74) := "11111111";
			tmp(54,75) := "11111111";
			tmp(54,76) := "11111111";
			tmp(54,77) := "11111111";
			tmp(54,78) := "11111111";
			tmp(54,79) := "11111111";
			tmp(54,80) := "11111111";
			tmp(55,1) := "11111111";
			tmp(55,2) := "11111110";
			tmp(55,3) := "11111110";
			tmp(55,4) := "11011101";
			tmp(55,5) := "00111001";
			tmp(55,6) := "00110001";
			tmp(55,7) := "01000100";
			tmp(55,8) := "01000110";
			tmp(55,9) := "01000000";
			tmp(55,10) := "01000110";
			tmp(55,11) := "01001101";
			tmp(55,12) := "10011101";
			tmp(55,13) := "10111100";
			tmp(55,14) := "11100001";
			tmp(55,15) := "11111001";
			tmp(55,16) := "11111111";
			tmp(55,17) := "11111100";
			tmp(55,18) := "11111111";
			tmp(55,19) := "11111101";
			tmp(55,20) := "11111111";
			tmp(55,21) := "11111110";
			tmp(55,22) := "11111100";
			tmp(55,23) := "11011011";
			tmp(55,24) := "01101110";
			tmp(55,25) := "10001100";
			tmp(55,26) := "11000010";
			tmp(55,27) := "11001100";
			tmp(55,28) := "10000101";
			tmp(55,29) := "01001000";
			tmp(55,30) := "01101110";
			tmp(55,31) := "01101010";
			tmp(55,32) := "01111001";
			tmp(55,33) := "01101010";
			tmp(55,34) := "10001011";
			tmp(55,35) := "10011101";
			tmp(55,36) := "10010111";
			tmp(55,37) := "10110010";
			tmp(55,38) := "10100010";
			tmp(55,39) := "10011110";
			tmp(55,40) := "10110010";
			tmp(55,41) := "10101100";
			tmp(55,42) := "10101100";
			tmp(55,43) := "10100011";
			tmp(55,44) := "10001111";
			tmp(55,45) := "10010010";
			tmp(55,46) := "10100001";
			tmp(55,47) := "10100001";
			tmp(55,48) := "10010101";
			tmp(55,49) := "10000111";
			tmp(55,50) := "01111111";
			tmp(55,51) := "10000110";
			tmp(55,52) := "01101110";
			tmp(55,53) := "10000110";
			tmp(55,54) := "01111010";
			tmp(55,55) := "01111100";
			tmp(55,56) := "10100100";
			tmp(55,57) := "10011110";
			tmp(55,58) := "01101111";
			tmp(55,59) := "10101101";
			tmp(55,60) := "11010001";
			tmp(55,61) := "11101000";
			tmp(55,62) := "11111000";
			tmp(55,63) := "11111111";
			tmp(55,64) := "11111111";
			tmp(55,65) := "11111011";
			tmp(55,66) := "11111111";
			tmp(55,67) := "11111110";
			tmp(55,68) := "11111111";
			tmp(55,69) := "11111111";
			tmp(55,70) := "11111111";
			tmp(55,71) := "11111110";
			tmp(55,72) := "11111110";
			tmp(55,73) := "11111111";
			tmp(55,74) := "11111111";
			tmp(55,75) := "11111111";
			tmp(55,76) := "11111111";
			tmp(55,77) := "11111111";
			tmp(55,78) := "11111111";
			tmp(55,79) := "11111111";
			tmp(55,80) := "11111111";
			tmp(56,1) := "11111100";
			tmp(56,2) := "11111111";
			tmp(56,3) := "11111111";
			tmp(56,4) := "11101010";
			tmp(56,5) := "11010101";
			tmp(56,6) := "11001000";
			tmp(56,7) := "11001110";
			tmp(56,8) := "11001111";
			tmp(56,9) := "11100010";
			tmp(56,10) := "11011110";
			tmp(56,11) := "11110001";
			tmp(56,12) := "11111000";
			tmp(56,13) := "11111100";
			tmp(56,14) := "11111110";
			tmp(56,15) := "11111110";
			tmp(56,16) := "11111110";
			tmp(56,17) := "11111111";
			tmp(56,18) := "11111010";
			tmp(56,19) := "11111100";
			tmp(56,20) := "11111111";
			tmp(56,21) := "11111111";
			tmp(56,22) := "11111101";
			tmp(56,23) := "10100010";
			tmp(56,24) := "01111101";
			tmp(56,25) := "10000010";
			tmp(56,26) := "10110001";
			tmp(56,27) := "11111010";
			tmp(56,28) := "10110001";
			tmp(56,29) := "01010100";
			tmp(56,30) := "01001110";
			tmp(56,31) := "01100000";
			tmp(56,32) := "01100000";
			tmp(56,33) := "01100110";
			tmp(56,34) := "01101100";
			tmp(56,35) := "01111000";
			tmp(56,36) := "10001010";
			tmp(56,37) := "10011010";
			tmp(56,38) := "10010111";
			tmp(56,39) := "10011010";
			tmp(56,40) := "10110011";
			tmp(56,41) := "10011110";
			tmp(56,42) := "10100101";
			tmp(56,43) := "10100101";
			tmp(56,44) := "10010010";
			tmp(56,45) := "10001000";
			tmp(56,46) := "10001100";
			tmp(56,47) := "10010001";
			tmp(56,48) := "10000011";
			tmp(56,49) := "10000011";
			tmp(56,50) := "01111001";
			tmp(56,51) := "01110111";
			tmp(56,52) := "10000011";
			tmp(56,53) := "10010010";
			tmp(56,54) := "10011110";
			tmp(56,55) := "10001111";
			tmp(56,56) := "10011110";
			tmp(56,57) := "10000100";
			tmp(56,58) := "10001010";
			tmp(56,59) := "11010100";
			tmp(56,60) := "11111011";
			tmp(56,61) := "11111100";
			tmp(56,62) := "11111010";
			tmp(56,63) := "11111111";
			tmp(56,64) := "11111110";
			tmp(56,65) := "11111111";
			tmp(56,66) := "11111111";
			tmp(56,67) := "11111111";
			tmp(56,68) := "11111110";
			tmp(56,69) := "11111111";
			tmp(56,70) := "11111111";
			tmp(56,71) := "11111111";
			tmp(56,72) := "11111111";
			tmp(56,73) := "11111111";
			tmp(56,74) := "11111111";
			tmp(56,75) := "11111111";
			tmp(56,76) := "11111111";
			tmp(56,77) := "11111111";
			tmp(56,78) := "11111111";
			tmp(56,79) := "11111111";
			tmp(56,80) := "11111111";
			tmp(57,1) := "11111111";
			tmp(57,2) := "11111111";
			tmp(57,3) := "11111111";
			tmp(57,4) := "11111111";
			tmp(57,5) := "11111111";
			tmp(57,6) := "11111111";
			tmp(57,7) := "11111111";
			tmp(57,8) := "11111111";
			tmp(57,9) := "11111111";
			tmp(57,10) := "11111111";
			tmp(57,11) := "11111111";
			tmp(57,12) := "11111111";
			tmp(57,13) := "11111111";
			tmp(57,14) := "11111111";
			tmp(57,15) := "11111111";
			tmp(57,16) := "11111111";
			tmp(57,17) := "11111111";
			tmp(57,18) := "11111011";
			tmp(57,19) := "11111111";
			tmp(57,20) := "11111110";
			tmp(57,21) := "11111111";
			tmp(57,22) := "11101011";
			tmp(57,23) := "01110101";
			tmp(57,24) := "01011110";
			tmp(57,25) := "10000111";
			tmp(57,26) := "01111101";
			tmp(57,27) := "11101111";
			tmp(57,28) := "11101111";
			tmp(57,29) := "01101111";
			tmp(57,30) := "00111001";
			tmp(57,31) := "01011110";
			tmp(57,32) := "01011010";
			tmp(57,33) := "01011011";
			tmp(57,34) := "01100101";
			tmp(57,35) := "01110101";
			tmp(57,36) := "01111111";
			tmp(57,37) := "10010001";
			tmp(57,38) := "01111100";
			tmp(57,39) := "10000110";
			tmp(57,40) := "10101000";
			tmp(57,41) := "10101110";
			tmp(57,42) := "10011110";
			tmp(57,43) := "10011111";
			tmp(57,44) := "10010000";
			tmp(57,45) := "10001110";
			tmp(57,46) := "10000000";
			tmp(57,47) := "01111101";
			tmp(57,48) := "01111111";
			tmp(57,49) := "10000000";
			tmp(57,50) := "01110001";
			tmp(57,51) := "01110010";
			tmp(57,52) := "10010000";
			tmp(57,53) := "10011100";
			tmp(57,54) := "10011011";
			tmp(57,55) := "10011100";
			tmp(57,56) := "10010011";
			tmp(57,57) := "10100000";
			tmp(57,58) := "11010100";
			tmp(57,59) := "11111010";
			tmp(57,60) := "11111100";
			tmp(57,61) := "11111011";
			tmp(57,62) := "11111110";
			tmp(57,63) := "11111111";
			tmp(57,64) := "11111111";
			tmp(57,65) := "11111111";
			tmp(57,66) := "11111111";
			tmp(57,67) := "11111111";
			tmp(57,68) := "11111111";
			tmp(57,69) := "11111111";
			tmp(57,70) := "11111111";
			tmp(57,71) := "11111111";
			tmp(57,72) := "11111111";
			tmp(57,73) := "11111111";
			tmp(57,74) := "11111111";
			tmp(57,75) := "11111111";
			tmp(57,76) := "11111111";
			tmp(57,77) := "11111111";
			tmp(57,78) := "11111111";
			tmp(57,79) := "11111111";
			tmp(57,80) := "11111111";
			tmp(58,1) := "11111111";
			tmp(58,2) := "11111111";
			tmp(58,3) := "11111111";
			tmp(58,4) := "11111111";
			tmp(58,5) := "11111111";
			tmp(58,6) := "11111111";
			tmp(58,7) := "11111111";
			tmp(58,8) := "11111111";
			tmp(58,9) := "11111111";
			tmp(58,10) := "11111111";
			tmp(58,11) := "11111111";
			tmp(58,12) := "11111111";
			tmp(58,13) := "11111111";
			tmp(58,14) := "11111111";
			tmp(58,15) := "11111111";
			tmp(58,16) := "11111111";
			tmp(58,17) := "11111111";
			tmp(58,18) := "11111010";
			tmp(58,19) := "11111111";
			tmp(58,20) := "11111111";
			tmp(58,21) := "11111110";
			tmp(58,22) := "11011011";
			tmp(58,23) := "01101011";
			tmp(58,24) := "01010110";
			tmp(58,25) := "01110011";
			tmp(58,26) := "01110011";
			tmp(58,27) := "10101110";
			tmp(58,28) := "11111110";
			tmp(58,29) := "10011010";
			tmp(58,30) := "01001000";
			tmp(58,31) := "01001011";
			tmp(58,32) := "01011111";
			tmp(58,33) := "01101000";
			tmp(58,34) := "01101001";
			tmp(58,35) := "01101110";
			tmp(58,36) := "01110010";
			tmp(58,37) := "01111001";
			tmp(58,38) := "01110101";
			tmp(58,39) := "01110110";
			tmp(58,40) := "10000100";
			tmp(58,41) := "10001110";
			tmp(58,42) := "10011011";
			tmp(58,43) := "10010001";
			tmp(58,44) := "10001000";
			tmp(58,45) := "10001010";
			tmp(58,46) := "01111100";
			tmp(58,47) := "01101101";
			tmp(58,48) := "10001000";
			tmp(58,49) := "10000101";
			tmp(58,50) := "10000010";
			tmp(58,51) := "10000110";
			tmp(58,52) := "10011111";
			tmp(58,53) := "10011001";
			tmp(58,54) := "10101000";
			tmp(58,55) := "01111001";
			tmp(58,56) := "10101110";
			tmp(58,57) := "11110110";
			tmp(58,58) := "11111110";
			tmp(58,59) := "11111110";
			tmp(58,60) := "11111110";
			tmp(58,61) := "11111111";
			tmp(58,62) := "11111111";
			tmp(58,63) := "11111111";
			tmp(58,64) := "11111111";
			tmp(58,65) := "11111111";
			tmp(58,66) := "11111111";
			tmp(58,67) := "11111111";
			tmp(58,68) := "11111111";
			tmp(58,69) := "11111111";
			tmp(58,70) := "11111111";
			tmp(58,71) := "11111111";
			tmp(58,72) := "11111111";
			tmp(58,73) := "11111111";
			tmp(58,74) := "11111111";
			tmp(58,75) := "11111111";
			tmp(58,76) := "11111111";
			tmp(58,77) := "11111111";
			tmp(58,78) := "11111111";
			tmp(58,79) := "11111111";
			tmp(58,80) := "11111111";
			tmp(59,1) := "11111111";
			tmp(59,2) := "11111111";
			tmp(59,3) := "11111111";
			tmp(59,4) := "11111111";
			tmp(59,5) := "11111111";
			tmp(59,6) := "11111111";
			tmp(59,7) := "11111111";
			tmp(59,8) := "11111111";
			tmp(59,9) := "11111111";
			tmp(59,10) := "11111111";
			tmp(59,11) := "11111111";
			tmp(59,12) := "11111111";
			tmp(59,13) := "11111111";
			tmp(59,14) := "11111111";
			tmp(59,15) := "11111111";
			tmp(59,16) := "11111111";
			tmp(59,17) := "11111111";
			tmp(59,18) := "11111100";
			tmp(59,19) := "11111111";
			tmp(59,20) := "11111111";
			tmp(59,21) := "11110111";
			tmp(59,22) := "11010000";
			tmp(59,23) := "00111100";
			tmp(59,24) := "01001011";
			tmp(59,25) := "01101000";
			tmp(59,26) := "01000111";
			tmp(59,27) := "10101110";
			tmp(59,28) := "11111011";
			tmp(59,29) := "11011001";
			tmp(59,30) := "00101011";
			tmp(59,31) := "00111101";
			tmp(59,32) := "01100010";
			tmp(59,33) := "01011111";
			tmp(59,34) := "01101011";
			tmp(59,35) := "01110010";
			tmp(59,36) := "01101110";
			tmp(59,37) := "01110111";
			tmp(59,38) := "10000100";
			tmp(59,39) := "10000001";
			tmp(59,40) := "01111100";
			tmp(59,41) := "10000011";
			tmp(59,42) := "10001101";
			tmp(59,43) := "10000011";
			tmp(59,44) := "10011010";
			tmp(59,45) := "10010010";
			tmp(59,46) := "10000101";
			tmp(59,47) := "01111110";
			tmp(59,48) := "10000001";
			tmp(59,49) := "10001000";
			tmp(59,50) := "10010000";
			tmp(59,51) := "10101011";
			tmp(59,52) := "10011101";
			tmp(59,53) := "10011011";
			tmp(59,54) := "10111000";
			tmp(59,55) := "11100000";
			tmp(59,56) := "11101100";
			tmp(59,57) := "11111011";
			tmp(59,58) := "11111011";
			tmp(59,59) := "11111011";
			tmp(59,60) := "11111110";
			tmp(59,61) := "11111111";
			tmp(59,62) := "11111111";
			tmp(59,63) := "11111101";
			tmp(59,64) := "11111000";
			tmp(59,65) := "11111111";
			tmp(59,66) := "11111111";
			tmp(59,67) := "11111111";
			tmp(59,68) := "11111111";
			tmp(59,69) := "11111111";
			tmp(59,70) := "11111111";
			tmp(59,71) := "11111111";
			tmp(59,72) := "11111111";
			tmp(59,73) := "11111111";
			tmp(59,74) := "11111111";
			tmp(59,75) := "11111111";
			tmp(59,76) := "11111111";
			tmp(59,77) := "11111111";
			tmp(59,78) := "11111111";
			tmp(59,79) := "11111111";
			tmp(59,80) := "11111111";
			tmp(60,1) := "11111111";
			tmp(60,2) := "11111111";
			tmp(60,3) := "11111111";
			tmp(60,4) := "11111111";
			tmp(60,5) := "11111111";
			tmp(60,6) := "11111111";
			tmp(60,7) := "11111111";
			tmp(60,8) := "11111111";
			tmp(60,9) := "11111111";
			tmp(60,10) := "11111111";
			tmp(60,11) := "11111111";
			tmp(60,12) := "11111111";
			tmp(60,13) := "11111111";
			tmp(60,14) := "11111111";
			tmp(60,15) := "11111111";
			tmp(60,16) := "11111111";
			tmp(60,17) := "11111111";
			tmp(60,18) := "11111110";
			tmp(60,19) := "11111111";
			tmp(60,20) := "11111110";
			tmp(60,21) := "11111000";
			tmp(60,22) := "10000100";
			tmp(60,23) := "00111010";
			tmp(60,24) := "00111101";
			tmp(60,25) := "01000101";
			tmp(60,26) := "01010000";
			tmp(60,27) := "01011000";
			tmp(60,28) := "11111111";
			tmp(60,29) := "11000100";
			tmp(60,30) := "00111100";
			tmp(60,31) := "00110111";
			tmp(60,32) := "01001101";
			tmp(60,33) := "01100101";
			tmp(60,34) := "01001101";
			tmp(60,35) := "01011011";
			tmp(60,36) := "01100011";
			tmp(60,37) := "01101101";
			tmp(60,38) := "01111110";
			tmp(60,39) := "10010101";
			tmp(60,40) := "10011100";
			tmp(60,41) := "10000111";
			tmp(60,42) := "10000011";
			tmp(60,43) := "10001001";
			tmp(60,44) := "10010111";
			tmp(60,45) := "10001111";
			tmp(60,46) := "10000100";
			tmp(60,47) := "10001010";
			tmp(60,48) := "10010111";
			tmp(60,49) := "01111111";
			tmp(60,50) := "10001001";
			tmp(60,51) := "10001110";
			tmp(60,52) := "10000001";
			tmp(60,53) := "10101001";
			tmp(60,54) := "11011000";
			tmp(60,55) := "11110101";
			tmp(60,56) := "11111011";
			tmp(60,57) := "11111111";
			tmp(60,58) := "11111111";
			tmp(60,59) := "11111111";
			tmp(60,60) := "11111111";
			tmp(60,61) := "11111111";
			tmp(60,62) := "11111111";
			tmp(60,63) := "11111110";
			tmp(60,64) := "11111011";
			tmp(60,65) := "11111111";
			tmp(60,66) := "11111111";
			tmp(60,67) := "11111111";
			tmp(60,68) := "11111111";
			tmp(60,69) := "11111111";
			tmp(60,70) := "11111111";
			tmp(60,71) := "11111111";
			tmp(60,72) := "11111111";
			tmp(60,73) := "11111111";
			tmp(60,74) := "11111111";
			tmp(60,75) := "11111111";
			tmp(60,76) := "11111111";
			tmp(60,77) := "11111111";
			tmp(60,78) := "11111111";
			tmp(60,79) := "11111111";
			tmp(60,80) := "11111111";
			tmp(61,1) := "11111111";
			tmp(61,2) := "11111111";
			tmp(61,3) := "11111111";
			tmp(61,4) := "11111111";
			tmp(61,5) := "11111111";
			tmp(61,6) := "11111111";
			tmp(61,7) := "11111111";
			tmp(61,8) := "11111111";
			tmp(61,9) := "11111111";
			tmp(61,10) := "11111111";
			tmp(61,11) := "11111111";
			tmp(61,12) := "11111111";
			tmp(61,13) := "11111111";
			tmp(61,14) := "11111111";
			tmp(61,15) := "11111111";
			tmp(61,16) := "11111111";
			tmp(61,17) := "11111111";
			tmp(61,18) := "11111111";
			tmp(61,19) := "11111111";
			tmp(61,20) := "11111111";
			tmp(61,21) := "11100001";
			tmp(61,22) := "01100101";
			tmp(61,23) := "00110101";
			tmp(61,24) := "00110100";
			tmp(61,25) := "00110111";
			tmp(61,26) := "00111010";
			tmp(61,27) := "01100111";
			tmp(61,28) := "11000110";
			tmp(61,29) := "11011001";
			tmp(61,30) := "00111101";
			tmp(61,31) := "01001000";
			tmp(61,32) := "01111111";
			tmp(61,33) := "01111001";
			tmp(61,34) := "01010000";
			tmp(61,35) := "01000010";
			tmp(61,36) := "01010111";
			tmp(61,37) := "01010001";
			tmp(61,38) := "01011111";
			tmp(61,39) := "01111011";
			tmp(61,40) := "10010001";
			tmp(61,41) := "10001101";
			tmp(61,42) := "10000101";
			tmp(61,43) := "10011100";
			tmp(61,44) := "11001001";
			tmp(61,45) := "10100011";
			tmp(61,46) := "10010100";
			tmp(61,47) := "10011001";
			tmp(61,48) := "10001111";
			tmp(61,49) := "10010010";
			tmp(61,50) := "10101011";
			tmp(61,51) := "10110100";
			tmp(61,52) := "11011010";
			tmp(61,53) := "11101010";
			tmp(61,54) := "11111010";
			tmp(61,55) := "11111100";
			tmp(61,56) := "11111111";
			tmp(61,57) := "11111111";
			tmp(61,58) := "11111110";
			tmp(61,59) := "11111101";
			tmp(61,60) := "11111110";
			tmp(61,61) := "11111111";
			tmp(61,62) := "11111111";
			tmp(61,63) := "11111111";
			tmp(61,64) := "11111111";
			tmp(61,65) := "11111111";
			tmp(61,66) := "11111111";
			tmp(61,67) := "11111111";
			tmp(61,68) := "11111111";
			tmp(61,69) := "11111111";
			tmp(61,70) := "11111111";
			tmp(61,71) := "11111111";
			tmp(61,72) := "11111111";
			tmp(61,73) := "11111111";
			tmp(61,74) := "11111111";
			tmp(61,75) := "11111111";
			tmp(61,76) := "11111111";
			tmp(61,77) := "11111111";
			tmp(61,78) := "11111111";
			tmp(61,79) := "11111111";
			tmp(61,80) := "11111111";
			tmp(62,1) := "11111111";
			tmp(62,2) := "11111111";
			tmp(62,3) := "11111111";
			tmp(62,4) := "11111111";
			tmp(62,5) := "11111111";
			tmp(62,6) := "11111111";
			tmp(62,7) := "11111111";
			tmp(62,8) := "11111111";
			tmp(62,9) := "11111111";
			tmp(62,10) := "11111111";
			tmp(62,11) := "11111111";
			tmp(62,12) := "11111111";
			tmp(62,13) := "11111111";
			tmp(62,14) := "11111111";
			tmp(62,15) := "11111111";
			tmp(62,16) := "11111111";
			tmp(62,17) := "11111111";
			tmp(62,18) := "11111110";
			tmp(62,19) := "11111111";
			tmp(62,20) := "11111111";
			tmp(62,21) := "11011001";
			tmp(62,22) := "01100001";
			tmp(62,23) := "00101011";
			tmp(62,24) := "00110100";
			tmp(62,25) := "00111100";
			tmp(62,26) := "00110100";
			tmp(62,27) := "00100011";
			tmp(62,28) := "10110101";
			tmp(62,29) := "10000001";
			tmp(62,30) := "01000000";
			tmp(62,31) := "01101110";
			tmp(62,32) := "10011010";
			tmp(62,33) := "10001001";
			tmp(62,34) := "01001111";
			tmp(62,35) := "00101110";
			tmp(62,36) := "01000111";
			tmp(62,37) := "01010110";
			tmp(62,38) := "01001000";
			tmp(62,39) := "10000101";
			tmp(62,40) := "11101101";
			tmp(62,41) := "11011110";
			tmp(62,42) := "11100010";
			tmp(62,43) := "11001011";
			tmp(62,44) := "10011000";
			tmp(62,45) := "10011010";
			tmp(62,46) := "10111011";
			tmp(62,47) := "11000111";
			tmp(62,48) := "10111001";
			tmp(62,49) := "11010100";
			tmp(62,50) := "11110010";
			tmp(62,51) := "11111100";
			tmp(62,52) := "11111100";
			tmp(62,53) := "11111100";
			tmp(62,54) := "11111111";
			tmp(62,55) := "11111111";
			tmp(62,56) := "11111101";
			tmp(62,57) := "11111100";
			tmp(62,58) := "11111011";
			tmp(62,59) := "11111110";
			tmp(62,60) := "11111111";
			tmp(62,61) := "11111111";
			tmp(62,62) := "11111111";
			tmp(62,63) := "11111111";
			tmp(62,64) := "11111111";
			tmp(62,65) := "11111111";
			tmp(62,66) := "11111111";
			tmp(62,67) := "11111111";
			tmp(62,68) := "11111111";
			tmp(62,69) := "11111111";
			tmp(62,70) := "11111111";
			tmp(62,71) := "11111111";
			tmp(62,72) := "11111111";
			tmp(62,73) := "11111111";
			tmp(62,74) := "11111111";
			tmp(62,75) := "11111111";
			tmp(62,76) := "11111111";
			tmp(62,77) := "11111111";
			tmp(62,78) := "11111111";
			tmp(62,79) := "11111111";
			tmp(62,80) := "11111111";
			tmp(63,1) := "11111111";
			tmp(63,2) := "11111111";
			tmp(63,3) := "11111111";
			tmp(63,4) := "11111111";
			tmp(63,5) := "11111111";
			tmp(63,6) := "11111111";
			tmp(63,7) := "11111111";
			tmp(63,8) := "11111111";
			tmp(63,9) := "11111111";
			tmp(63,10) := "11111111";
			tmp(63,11) := "11111111";
			tmp(63,12) := "11111111";
			tmp(63,13) := "11111111";
			tmp(63,14) := "11111111";
			tmp(63,15) := "11111111";
			tmp(63,16) := "11111111";
			tmp(63,17) := "11111110";
			tmp(63,18) := "11111111";
			tmp(63,19) := "11111110";
			tmp(63,20) := "11111100";
			tmp(63,21) := "11011001";
			tmp(63,22) := "00101100";
			tmp(63,23) := "00111001";
			tmp(63,24) := "00101100";
			tmp(63,25) := "00101100";
			tmp(63,26) := "00110111";
			tmp(63,27) := "00111001";
			tmp(63,28) := "01010000";
			tmp(63,29) := "01100101";
			tmp(63,30) := "01010011";
			tmp(63,31) := "01011101";
			tmp(63,32) := "10001011";
			tmp(63,33) := "01111111";
			tmp(63,34) := "01001101";
			tmp(63,35) := "00111001";
			tmp(63,36) := "00110110";
			tmp(63,37) := "01010110";
			tmp(63,38) := "00111100";
			tmp(63,39) := "01101011";
			tmp(63,40) := "11100011";
			tmp(63,41) := "11111111";
			tmp(63,42) := "11111111";
			tmp(63,43) := "11111101";
			tmp(63,44) := "11110111";
			tmp(63,45) := "11111010";
			tmp(63,46) := "11111011";
			tmp(63,47) := "11111111";
			tmp(63,48) := "11111111";
			tmp(63,49) := "11111111";
			tmp(63,50) := "11111011";
			tmp(63,51) := "11111010";
			tmp(63,52) := "11111111";
			tmp(63,53) := "11111110";
			tmp(63,54) := "11111100";
			tmp(63,55) := "11111111";
			tmp(63,56) := "11111111";
			tmp(63,57) := "11111111";
			tmp(63,58) := "11111111";
			tmp(63,59) := "11111111";
			tmp(63,60) := "11111101";
			tmp(63,61) := "11111110";
			tmp(63,62) := "11111110";
			tmp(63,63) := "11111100";
			tmp(63,64) := "11111100";
			tmp(63,65) := "11111111";
			tmp(63,66) := "11111111";
			tmp(63,67) := "11111111";
			tmp(63,68) := "11111111";
			tmp(63,69) := "11111111";
			tmp(63,70) := "11111111";
			tmp(63,71) := "11111111";
			tmp(63,72) := "11111111";
			tmp(63,73) := "11111111";
			tmp(63,74) := "11111111";
			tmp(63,75) := "11111111";
			tmp(63,76) := "11111111";
			tmp(63,77) := "11111111";
			tmp(63,78) := "11111111";
			tmp(63,79) := "11111111";
			tmp(63,80) := "11111111";
			tmp(64,1) := "11111111";
			tmp(64,2) := "11111111";
			tmp(64,3) := "11111111";
			tmp(64,4) := "11111111";
			tmp(64,5) := "11111111";
			tmp(64,6) := "11111111";
			tmp(64,7) := "11111111";
			tmp(64,8) := "11111111";
			tmp(64,9) := "11111111";
			tmp(64,10) := "11111111";
			tmp(64,11) := "11111111";
			tmp(64,12) := "11111111";
			tmp(64,13) := "11111111";
			tmp(64,14) := "11111111";
			tmp(64,15) := "11111111";
			tmp(64,16) := "11111111";
			tmp(64,17) := "11111100";
			tmp(64,18) := "11111111";
			tmp(64,19) := "11111100";
			tmp(64,20) := "11111111";
			tmp(64,21) := "10110101";
			tmp(64,22) := "01001100";
			tmp(64,23) := "00111000";
			tmp(64,24) := "00110001";
			tmp(64,25) := "00101101";
			tmp(64,26) := "00101001";
			tmp(64,27) := "00110110";
			tmp(64,28) := "10011011";
			tmp(64,29) := "10000001";
			tmp(64,30) := "01000110";
			tmp(64,31) := "01000110";
			tmp(64,32) := "01010001";
			tmp(64,33) := "10000001";
			tmp(64,34) := "01011011";
			tmp(64,35) := "00101101";
			tmp(64,36) := "00100011";
			tmp(64,37) := "00111101";
			tmp(64,38) := "01010100";
			tmp(64,39) := "01010111";
			tmp(64,40) := "11011111";
			tmp(64,41) := "11111011";
			tmp(64,42) := "11111101";
			tmp(64,43) := "11111111";
			tmp(64,44) := "11111111";
			tmp(64,45) := "11111011";
			tmp(64,46) := "11111110";
			tmp(64,47) := "11111111";
			tmp(64,48) := "11111111";
			tmp(64,49) := "11111111";
			tmp(64,50) := "11111111";
			tmp(64,51) := "11111111";
			tmp(64,52) := "11111101";
			tmp(64,53) := "11111111";
			tmp(64,54) := "11111111";
			tmp(64,55) := "11111100";
			tmp(64,56) := "11111110";
			tmp(64,57) := "11111111";
			tmp(64,58) := "11111111";
			tmp(64,59) := "11111111";
			tmp(64,60) := "11111111";
			tmp(64,61) := "11111111";
			tmp(64,62) := "11111111";
			tmp(64,63) := "11111111";
			tmp(64,64) := "11111111";
			tmp(64,65) := "11111111";
			tmp(64,66) := "11111111";
			tmp(64,67) := "11111111";
			tmp(64,68) := "11111111";
			tmp(64,69) := "11111111";
			tmp(64,70) := "11111111";
			tmp(64,71) := "11111111";
			tmp(64,72) := "11111111";
			tmp(64,73) := "11111111";
			tmp(64,74) := "11111111";
			tmp(64,75) := "11111111";
			tmp(64,76) := "11111111";
			tmp(64,77) := "11111111";
			tmp(64,78) := "11111111";
			tmp(64,79) := "11111111";
			tmp(64,80) := "11111111";
			tmp(65,1) := "11111111";
			tmp(65,2) := "11111111";
			tmp(65,3) := "11111111";
			tmp(65,4) := "11111111";
			tmp(65,5) := "11111111";
			tmp(65,6) := "11111111";
			tmp(65,7) := "11111111";
			tmp(65,8) := "11111111";
			tmp(65,9) := "11111111";
			tmp(65,10) := "11111111";
			tmp(65,11) := "11111111";
			tmp(65,12) := "11111111";
			tmp(65,13) := "11111111";
			tmp(65,14) := "11111111";
			tmp(65,15) := "11111111";
			tmp(65,16) := "11111111";
			tmp(65,17) := "11111111";
			tmp(65,18) := "11111011";
			tmp(65,19) := "11111110";
			tmp(65,20) := "11111111";
			tmp(65,21) := "11011000";
			tmp(65,22) := "00111011";
			tmp(65,23) := "01000111";
			tmp(65,24) := "00111100";
			tmp(65,25) := "00110110";
			tmp(65,26) := "00101000";
			tmp(65,27) := "01001000";
			tmp(65,28) := "10000111";
			tmp(65,29) := "10001110";
			tmp(65,30) := "01001110";
			tmp(65,31) := "00111110";
			tmp(65,32) := "00111101";
			tmp(65,33) := "01101110";
			tmp(65,34) := "01111011";
			tmp(65,35) := "00111010";
			tmp(65,36) := "00101100";
			tmp(65,37) := "00101110";
			tmp(65,38) := "01001001";
			tmp(65,39) := "01011101";
			tmp(65,40) := "11010000";
			tmp(65,41) := "11111110";
			tmp(65,42) := "11111110";
			tmp(65,43) := "11111111";
			tmp(65,44) := "11111110";
			tmp(65,45) := "11111111";
			tmp(65,46) := "11111111";
			tmp(65,47) := "11111111";
			tmp(65,48) := "11111111";
			tmp(65,49) := "11111111";
			tmp(65,50) := "11111111";
			tmp(65,51) := "11111111";
			tmp(65,52) := "11111111";
			tmp(65,53) := "11111111";
			tmp(65,54) := "11111111";
			tmp(65,55) := "11111111";
			tmp(65,56) := "11111111";
			tmp(65,57) := "11111111";
			tmp(65,58) := "11111111";
			tmp(65,59) := "11111111";
			tmp(65,60) := "11111111";
			tmp(65,61) := "11111111";
			tmp(65,62) := "11111111";
			tmp(65,63) := "11111111";
			tmp(65,64) := "11111111";
			tmp(65,65) := "11111111";
			tmp(65,66) := "11111111";
			tmp(65,67) := "11111111";
			tmp(65,68) := "11111111";
			tmp(65,69) := "11111111";
			tmp(65,70) := "11111111";
			tmp(65,71) := "11111111";
			tmp(65,72) := "11111111";
			tmp(65,73) := "11111111";
			tmp(65,74) := "11111111";
			tmp(65,75) := "11111111";
			tmp(65,76) := "11111111";
			tmp(65,77) := "11111111";
			tmp(65,78) := "11111111";
			tmp(65,79) := "11111111";
			tmp(65,80) := "11111111";
			tmp(66,1) := "11111111";
			tmp(66,2) := "11111111";
			tmp(66,3) := "11111111";
			tmp(66,4) := "11111111";
			tmp(66,5) := "11111111";
			tmp(66,6) := "11111111";
			tmp(66,7) := "11111111";
			tmp(66,8) := "11111111";
			tmp(66,9) := "11111111";
			tmp(66,10) := "11111111";
			tmp(66,11) := "11111111";
			tmp(66,12) := "11111111";
			tmp(66,13) := "11111111";
			tmp(66,14) := "11111111";
			tmp(66,15) := "11111111";
			tmp(66,16) := "11111111";
			tmp(66,17) := "11111111";
			tmp(66,18) := "11111100";
			tmp(66,19) := "11111111";
			tmp(66,20) := "11111111";
			tmp(66,21) := "11000011";
			tmp(66,22) := "01100101";
			tmp(66,23) := "01000101";
			tmp(66,24) := "01000001";
			tmp(66,25) := "00111100";
			tmp(66,26) := "00101111";
			tmp(66,27) := "00101110";
			tmp(66,28) := "01100011";
			tmp(66,29) := "01010101";
			tmp(66,30) := "00111001";
			tmp(66,31) := "01000101";
			tmp(66,32) := "00111100";
			tmp(66,33) := "00110011";
			tmp(66,34) := "01111110";
			tmp(66,35) := "01100010";
			tmp(66,36) := "00111100";
			tmp(66,37) := "01000011";
			tmp(66,38) := "00101001";
			tmp(66,39) := "01001101";
			tmp(66,40) := "11011111";
			tmp(66,41) := "11111100";
			tmp(66,42) := "11111111";
			tmp(66,43) := "11111111";
			tmp(66,44) := "11111110";
			tmp(66,45) := "11111100";
			tmp(66,46) := "11111111";
			tmp(66,47) := "11111111";
			tmp(66,48) := "11111110";
			tmp(66,49) := "11111111";
			tmp(66,50) := "11111111";
			tmp(66,51) := "11111111";
			tmp(66,52) := "11111111";
			tmp(66,53) := "11111111";
			tmp(66,54) := "11111111";
			tmp(66,55) := "11111111";
			tmp(66,56) := "11111111";
			tmp(66,57) := "11111111";
			tmp(66,58) := "11111111";
			tmp(66,59) := "11111111";
			tmp(66,60) := "11111111";
			tmp(66,61) := "11111111";
			tmp(66,62) := "11111111";
			tmp(66,63) := "11111111";
			tmp(66,64) := "11111111";
			tmp(66,65) := "11111111";
			tmp(66,66) := "11111111";
			tmp(66,67) := "11111111";
			tmp(66,68) := "11111111";
			tmp(66,69) := "11111111";
			tmp(66,70) := "11111111";
			tmp(66,71) := "11111111";
			tmp(66,72) := "11111111";
			tmp(66,73) := "11111111";
			tmp(66,74) := "11111111";
			tmp(66,75) := "11111111";
			tmp(66,76) := "11111111";
			tmp(66,77) := "11111111";
			tmp(66,78) := "11111111";
			tmp(66,79) := "11111111";
			tmp(66,80) := "11111111";
			tmp(67,1) := "11111111";
			tmp(67,2) := "11111111";
			tmp(67,3) := "11111111";
			tmp(67,4) := "11111111";
			tmp(67,5) := "11111111";
			tmp(67,6) := "11111111";
			tmp(67,7) := "11111111";
			tmp(67,8) := "11111111";
			tmp(67,9) := "11111111";
			tmp(67,10) := "11111111";
			tmp(67,11) := "11111111";
			tmp(67,12) := "11111111";
			tmp(67,13) := "11111111";
			tmp(67,14) := "11111111";
			tmp(67,15) := "11111111";
			tmp(67,16) := "11111111";
			tmp(67,17) := "11111111";
			tmp(67,18) := "11111100";
			tmp(67,19) := "11111110";
			tmp(67,20) := "11111111";
			tmp(67,21) := "11110000";
			tmp(67,22) := "01100001";
			tmp(67,23) := "01010100";
			tmp(67,24) := "01000100";
			tmp(67,25) := "00111101";
			tmp(67,26) := "00110100";
			tmp(67,27) := "00111000";
			tmp(67,28) := "01100011";
			tmp(67,29) := "01000111";
			tmp(67,30) := "01000001";
			tmp(67,31) := "01000100";
			tmp(67,32) := "00111011";
			tmp(67,33) := "00110101";
			tmp(67,34) := "01001011";
			tmp(67,35) := "01110101";
			tmp(67,36) := "01000110";
			tmp(67,37) := "01010010";
			tmp(67,38) := "01000010";
			tmp(67,39) := "00110010";
			tmp(67,40) := "10110001";
			tmp(67,41) := "11111110";
			tmp(67,42) := "11111111";
			tmp(67,43) := "11111111";
			tmp(67,44) := "11111101";
			tmp(67,45) := "11111110";
			tmp(67,46) := "11111100";
			tmp(67,47) := "11111111";
			tmp(67,48) := "11111011";
			tmp(67,49) := "11111111";
			tmp(67,50) := "11111111";
			tmp(67,51) := "11111111";
			tmp(67,52) := "11111111";
			tmp(67,53) := "11111111";
			tmp(67,54) := "11111111";
			tmp(67,55) := "11111111";
			tmp(67,56) := "11111111";
			tmp(67,57) := "11111111";
			tmp(67,58) := "11111111";
			tmp(67,59) := "11111111";
			tmp(67,60) := "11111111";
			tmp(67,61) := "11111111";
			tmp(67,62) := "11111111";
			tmp(67,63) := "11111111";
			tmp(67,64) := "11111111";
			tmp(67,65) := "11111111";
			tmp(67,66) := "11111111";
			tmp(67,67) := "11111111";
			tmp(67,68) := "11111111";
			tmp(67,69) := "11111111";
			tmp(67,70) := "11111111";
			tmp(67,71) := "11111111";
			tmp(67,72) := "11111111";
			tmp(67,73) := "11111111";
			tmp(67,74) := "11111111";
			tmp(67,75) := "11111111";
			tmp(67,76) := "11111111";
			tmp(67,77) := "11111111";
			tmp(67,78) := "11111111";
			tmp(67,79) := "11111111";
			tmp(67,80) := "11111111";
			tmp(68,1) := "11111111";
			tmp(68,2) := "11111111";
			tmp(68,3) := "11111111";
			tmp(68,4) := "11111111";
			tmp(68,5) := "11111111";
			tmp(68,6) := "11111111";
			tmp(68,7) := "11111111";
			tmp(68,8) := "11111111";
			tmp(68,9) := "11111111";
			tmp(68,10) := "11111111";
			tmp(68,11) := "11111111";
			tmp(68,12) := "11111111";
			tmp(68,13) := "11111111";
			tmp(68,14) := "11111111";
			tmp(68,15) := "11111111";
			tmp(68,16) := "11111111";
			tmp(68,17) := "11111101";
			tmp(68,18) := "11111111";
			tmp(68,19) := "11111110";
			tmp(68,20) := "11111101";
			tmp(68,21) := "11110101";
			tmp(68,22) := "10100011";
			tmp(68,23) := "01000111";
			tmp(68,24) := "01000000";
			tmp(68,25) := "01000010";
			tmp(68,26) := "00110110";
			tmp(68,27) := "01001001";
			tmp(68,28) := "01011110";
			tmp(68,29) := "01001111";
			tmp(68,30) := "00110111";
			tmp(68,31) := "01000001";
			tmp(68,32) := "01000011";
			tmp(68,33) := "00110100";
			tmp(68,34) := "01001010";
			tmp(68,35) := "01100000";
			tmp(68,36) := "01011110";
			tmp(68,37) := "01010111";
			tmp(68,38) := "01001001";
			tmp(68,39) := "01000000";
			tmp(68,40) := "01011000";
			tmp(68,41) := "11101011";
			tmp(68,42) := "11111111";
			tmp(68,43) := "11111111";
			tmp(68,44) := "11111111";
			tmp(68,45) := "11111011";
			tmp(68,46) := "11111111";
			tmp(68,47) := "11111111";
			tmp(68,48) := "11111100";
			tmp(68,49) := "11111111";
			tmp(68,50) := "11111111";
			tmp(68,51) := "11111111";
			tmp(68,52) := "11111111";
			tmp(68,53) := "11111111";
			tmp(68,54) := "11111111";
			tmp(68,55) := "11111111";
			tmp(68,56) := "11111111";
			tmp(68,57) := "11111111";
			tmp(68,58) := "11111111";
			tmp(68,59) := "11111111";
			tmp(68,60) := "11111111";
			tmp(68,61) := "11111111";
			tmp(68,62) := "11111111";
			tmp(68,63) := "11111111";
			tmp(68,64) := "11111111";
			tmp(68,65) := "11111111";
			tmp(68,66) := "11111111";
			tmp(68,67) := "11111111";
			tmp(68,68) := "11111111";
			tmp(68,69) := "11111111";
			tmp(68,70) := "11111111";
			tmp(68,71) := "11111111";
			tmp(68,72) := "11111111";
			tmp(68,73) := "11111111";
			tmp(68,74) := "11111111";
			tmp(68,75) := "11111111";
			tmp(68,76) := "11111111";
			tmp(68,77) := "11111111";
			tmp(68,78) := "11111111";
			tmp(68,79) := "11111111";
			tmp(68,80) := "11111111";
			tmp(69,1) := "11111111";
			tmp(69,2) := "11111111";
			tmp(69,3) := "11111111";
			tmp(69,4) := "11111111";
			tmp(69,5) := "11111111";
			tmp(69,6) := "11111111";
			tmp(69,7) := "11111111";
			tmp(69,8) := "11111111";
			tmp(69,9) := "11111111";
			tmp(69,10) := "11111111";
			tmp(69,11) := "11111111";
			tmp(69,12) := "11111111";
			tmp(69,13) := "11111111";
			tmp(69,14) := "11111111";
			tmp(69,15) := "11111111";
			tmp(69,16) := "11111111";
			tmp(69,17) := "11111110";
			tmp(69,18) := "11111110";
			tmp(69,19) := "11111110";
			tmp(69,20) := "11111111";
			tmp(69,21) := "11110110";
			tmp(69,22) := "10110111";
			tmp(69,23) := "01011000";
			tmp(69,24) := "00111100";
			tmp(69,25) := "01000100";
			tmp(69,26) := "00111011";
			tmp(69,27) := "01010111";
			tmp(69,28) := "10010011";
			tmp(69,29) := "00111000";
			tmp(69,30) := "00110011";
			tmp(69,31) := "00111110";
			tmp(69,32) := "01000000";
			tmp(69,33) := "00110110";
			tmp(69,34) := "00111001";
			tmp(69,35) := "01110101";
			tmp(69,36) := "01101011";
			tmp(69,37) := "01000111";
			tmp(69,38) := "01101011";
			tmp(69,39) := "01100111";
			tmp(69,40) := "01101011";
			tmp(69,41) := "10110100";
			tmp(69,42) := "11111011";
			tmp(69,43) := "11111100";
			tmp(69,44) := "11111111";
			tmp(69,45) := "11111111";
			tmp(69,46) := "11111111";
			tmp(69,47) := "11111111";
			tmp(69,48) := "11111110";
			tmp(69,49) := "11111111";
			tmp(69,50) := "11111111";
			tmp(69,51) := "11111111";
			tmp(69,52) := "11111111";
			tmp(69,53) := "11111111";
			tmp(69,54) := "11111111";
			tmp(69,55) := "11111111";
			tmp(69,56) := "11111111";
			tmp(69,57) := "11111111";
			tmp(69,58) := "11111111";
			tmp(69,59) := "11111111";
			tmp(69,60) := "11111111";
			tmp(69,61) := "11111111";
			tmp(69,62) := "11111111";
			tmp(69,63) := "11111111";
			tmp(69,64) := "11111111";
			tmp(69,65) := "11111111";
			tmp(69,66) := "11111111";
			tmp(69,67) := "11111111";
			tmp(69,68) := "11111111";
			tmp(69,69) := "11111111";
			tmp(69,70) := "11111111";
			tmp(69,71) := "11111111";
			tmp(69,72) := "11111111";
			tmp(69,73) := "11111111";
			tmp(69,74) := "11111111";
			tmp(69,75) := "11111111";
			tmp(69,76) := "11111111";
			tmp(69,77) := "11111111";
			tmp(69,78) := "11111111";
			tmp(69,79) := "11111111";
			tmp(69,80) := "11111111";
			tmp(70,1) := "11111111";
			tmp(70,2) := "11111111";
			tmp(70,3) := "11111111";
			tmp(70,4) := "11111111";
			tmp(70,5) := "11111111";
			tmp(70,6) := "11111111";
			tmp(70,7) := "11111111";
			tmp(70,8) := "11111111";
			tmp(70,9) := "11111111";
			tmp(70,10) := "11111111";
			tmp(70,11) := "11111111";
			tmp(70,12) := "11111111";
			tmp(70,13) := "11111111";
			tmp(70,14) := "11111111";
			tmp(70,15) := "11111111";
			tmp(70,16) := "11111111";
			tmp(70,17) := "11111110";
			tmp(70,18) := "11111111";
			tmp(70,19) := "11111101";
			tmp(70,20) := "11111111";
			tmp(70,21) := "11111111";
			tmp(70,22) := "11011110";
			tmp(70,23) := "01011000";
			tmp(70,24) := "01000000";
			tmp(70,25) := "01000000";
			tmp(70,26) := "00101111";
			tmp(70,27) := "10110011";
			tmp(70,28) := "10011001";
			tmp(70,29) := "01000001";
			tmp(70,30) := "00110000";
			tmp(70,31) := "00111101";
			tmp(70,32) := "00111110";
			tmp(70,33) := "00110101";
			tmp(70,34) := "00111001";
			tmp(70,35) := "01100100";
			tmp(70,36) := "01110010";
			tmp(70,37) := "01100110";
			tmp(70,38) := "10000011";
			tmp(70,39) := "11110101";
			tmp(70,40) := "10010010";
			tmp(70,41) := "10100111";
			tmp(70,42) := "11110010";
			tmp(70,43) := "11111111";
			tmp(70,44) := "11111111";
			tmp(70,45) := "11111111";
			tmp(70,46) := "11111111";
			tmp(70,47) := "11111110";
			tmp(70,48) := "11111111";
			tmp(70,49) := "11111111";
			tmp(70,50) := "11111111";
			tmp(70,51) := "11111111";
			tmp(70,52) := "11111111";
			tmp(70,53) := "11111111";
			tmp(70,54) := "11111111";
			tmp(70,55) := "11111111";
			tmp(70,56) := "11111111";
			tmp(70,57) := "11111111";
			tmp(70,58) := "11111111";
			tmp(70,59) := "11111111";
			tmp(70,60) := "11111111";
			tmp(70,61) := "11111111";
			tmp(70,62) := "11111111";
			tmp(70,63) := "11111111";
			tmp(70,64) := "11111111";
			tmp(70,65) := "11111111";
			tmp(70,66) := "11111111";
			tmp(70,67) := "11111111";
			tmp(70,68) := "11111111";
			tmp(70,69) := "11111111";
			tmp(70,70) := "11111111";
			tmp(70,71) := "11111111";
			tmp(70,72) := "11111111";
			tmp(70,73) := "11111111";
			tmp(70,74) := "11111111";
			tmp(70,75) := "11111111";
			tmp(70,76) := "11111111";
			tmp(70,77) := "11111111";
			tmp(70,78) := "11111111";
			tmp(70,79) := "11111111";
			tmp(70,80) := "11111111";
			tmp(71,1) := "11111111";
			tmp(71,2) := "11111111";
			tmp(71,3) := "11111111";
			tmp(71,4) := "11111111";
			tmp(71,5) := "11111111";
			tmp(71,6) := "11111111";
			tmp(71,7) := "11111111";
			tmp(71,8) := "11111111";
			tmp(71,9) := "11111111";
			tmp(71,10) := "11111111";
			tmp(71,11) := "11111111";
			tmp(71,12) := "11111111";
			tmp(71,13) := "11111111";
			tmp(71,14) := "11111111";
			tmp(71,15) := "11111111";
			tmp(71,16) := "11111111";
			tmp(71,17) := "11111111";
			tmp(71,18) := "11111110";
			tmp(71,19) := "11111111";
			tmp(71,20) := "11111110";
			tmp(71,21) := "11111111";
			tmp(71,22) := "11110110";
			tmp(71,23) := "10001111";
			tmp(71,24) := "01000101";
			tmp(71,25) := "00111101";
			tmp(71,26) := "01100110";
			tmp(71,27) := "11000011";
			tmp(71,28) := "11100110";
			tmp(71,29) := "01001101";
			tmp(71,30) := "00101011";
			tmp(71,31) := "00111000";
			tmp(71,32) := "00111100";
			tmp(71,33) := "00110101";
			tmp(71,34) := "00110101";
			tmp(71,35) := "01101101";
			tmp(71,36) := "01110000";
			tmp(71,37) := "10010001";
			tmp(71,38) := "11110011";
			tmp(71,39) := "11111101";
			tmp(71,40) := "11101100";
			tmp(71,41) := "10000010";
			tmp(71,42) := "11110111";
			tmp(71,43) := "11111111";
			tmp(71,44) := "11111111";
			tmp(71,45) := "11111111";
			tmp(71,46) := "11111111";
			tmp(71,47) := "11111111";
			tmp(71,48) := "11111101";
			tmp(71,49) := "11111111";
			tmp(71,50) := "11111111";
			tmp(71,51) := "11111111";
			tmp(71,52) := "11111111";
			tmp(71,53) := "11111111";
			tmp(71,54) := "11111111";
			tmp(71,55) := "11111111";
			tmp(71,56) := "11111111";
			tmp(71,57) := "11111111";
			tmp(71,58) := "11111111";
			tmp(71,59) := "11111111";
			tmp(71,60) := "11111111";
			tmp(71,61) := "11111111";
			tmp(71,62) := "11111111";
			tmp(71,63) := "11111111";
			tmp(71,64) := "11111111";
			tmp(71,65) := "11111111";
			tmp(71,66) := "11111111";
			tmp(71,67) := "11111111";
			tmp(71,68) := "11111111";
			tmp(71,69) := "11111111";
			tmp(71,70) := "11111111";
			tmp(71,71) := "11111111";
			tmp(71,72) := "11111111";
			tmp(71,73) := "11111111";
			tmp(71,74) := "11111111";
			tmp(71,75) := "11111111";
			tmp(71,76) := "11111111";
			tmp(71,77) := "11111111";
			tmp(71,78) := "11111111";
			tmp(71,79) := "11111111";
			tmp(71,80) := "11111111";
			tmp(72,1) := "11111111";
			tmp(72,2) := "11111111";
			tmp(72,3) := "11111111";
			tmp(72,4) := "11111111";
			tmp(72,5) := "11111111";
			tmp(72,6) := "11111111";
			tmp(72,7) := "11111111";
			tmp(72,8) := "11111111";
			tmp(72,9) := "11111111";
			tmp(72,10) := "11111111";
			tmp(72,11) := "11111111";
			tmp(72,12) := "11111111";
			tmp(72,13) := "11111111";
			tmp(72,14) := "11111111";
			tmp(72,15) := "11111111";
			tmp(72,16) := "11111111";
			tmp(72,17) := "11111111";
			tmp(72,18) := "11111011";
			tmp(72,19) := "11111111";
			tmp(72,20) := "11111111";
			tmp(72,21) := "11111110";
			tmp(72,22) := "11111101";
			tmp(72,23) := "11100000";
			tmp(72,24) := "01011011";
			tmp(72,25) := "00111110";
			tmp(72,26) := "01101001";
			tmp(72,27) := "11101110";
			tmp(72,28) := "11100110";
			tmp(72,29) := "01110101";
			tmp(72,30) := "00100011";
			tmp(72,31) := "00101100";
			tmp(72,32) := "00101111";
			tmp(72,33) := "00110111";
			tmp(72,34) := "10000001";
			tmp(72,35) := "10010111";
			tmp(72,36) := "10010101";
			tmp(72,37) := "11011100";
			tmp(72,38) := "11111110";
			tmp(72,39) := "11111111";
			tmp(72,40) := "11110101";
			tmp(72,41) := "11010100";
			tmp(72,42) := "11101000";
			tmp(72,43) := "11111111";
			tmp(72,44) := "11111111";
			tmp(72,45) := "11111101";
			tmp(72,46) := "11111110";
			tmp(72,47) := "11111101";
			tmp(72,48) := "11111100";
			tmp(72,49) := "11111111";
			tmp(72,50) := "11111111";
			tmp(72,51) := "11111111";
			tmp(72,52) := "11111111";
			tmp(72,53) := "11111111";
			tmp(72,54) := "11111111";
			tmp(72,55) := "11111111";
			tmp(72,56) := "11111111";
			tmp(72,57) := "11111111";
			tmp(72,58) := "11111111";
			tmp(72,59) := "11111111";
			tmp(72,60) := "11111111";
			tmp(72,61) := "11111111";
			tmp(72,62) := "11111111";
			tmp(72,63) := "11111111";
			tmp(72,64) := "11111111";
			tmp(72,65) := "11111111";
			tmp(72,66) := "11111111";
			tmp(72,67) := "11111111";
			tmp(72,68) := "11111111";
			tmp(72,69) := "11111111";
			tmp(72,70) := "11111111";
			tmp(72,71) := "11111111";
			tmp(72,72) := "11111111";
			tmp(72,73) := "11111111";
			tmp(72,74) := "11111111";
			tmp(72,75) := "11111111";
			tmp(72,76) := "11111111";
			tmp(72,77) := "11111111";
			tmp(72,78) := "11111111";
			tmp(72,79) := "11111111";
			tmp(72,80) := "11111111";
			tmp(73,1) := "11111111";
			tmp(73,2) := "11111111";
			tmp(73,3) := "11111111";
			tmp(73,4) := "11111111";
			tmp(73,5) := "11111111";
			tmp(73,6) := "11111111";
			tmp(73,7) := "11111111";
			tmp(73,8) := "11111111";
			tmp(73,9) := "11111111";
			tmp(73,10) := "11111111";
			tmp(73,11) := "11111111";
			tmp(73,12) := "11111111";
			tmp(73,13) := "11111111";
			tmp(73,14) := "11111111";
			tmp(73,15) := "11111111";
			tmp(73,16) := "11111111";
			tmp(73,17) := "11111111";
			tmp(73,18) := "11111111";
			tmp(73,19) := "11111111";
			tmp(73,20) := "11111111";
			tmp(73,21) := "11111101";
			tmp(73,22) := "11111111";
			tmp(73,23) := "11111101";
			tmp(73,24) := "11100011";
			tmp(73,25) := "01011011";
			tmp(73,26) := "10001010";
			tmp(73,27) := "11111000";
			tmp(73,28) := "11111011";
			tmp(73,29) := "11001111";
			tmp(73,30) := "10100010";
			tmp(73,31) := "10000011";
			tmp(73,32) := "10011100";
			tmp(73,33) := "11001010";
			tmp(73,34) := "11100011";
			tmp(73,35) := "11100100";
			tmp(73,36) := "10001111";
			tmp(73,37) := "11101101";
			tmp(73,38) := "11111111";
			tmp(73,39) := "11111111";
			tmp(73,40) := "11111010";
			tmp(73,41) := "11011110";
			tmp(73,42) := "11110110";
			tmp(73,43) := "11111110";
			tmp(73,44) := "11111101";
			tmp(73,45) := "11111111";
			tmp(73,46) := "11111111";
			tmp(73,47) := "11111110";
			tmp(73,48) := "11111111";
			tmp(73,49) := "11111111";
			tmp(73,50) := "11111111";
			tmp(73,51) := "11111111";
			tmp(73,52) := "11111111";
			tmp(73,53) := "11111111";
			tmp(73,54) := "11111111";
			tmp(73,55) := "11111111";
			tmp(73,56) := "11111111";
			tmp(73,57) := "11111111";
			tmp(73,58) := "11111111";
			tmp(73,59) := "11111111";
			tmp(73,60) := "11111111";
			tmp(73,61) := "11111111";
			tmp(73,62) := "11111111";
			tmp(73,63) := "11111111";
			tmp(73,64) := "11111111";
			tmp(73,65) := "11111111";
			tmp(73,66) := "11111111";
			tmp(73,67) := "11111111";
			tmp(73,68) := "11111111";
			tmp(73,69) := "11111111";
			tmp(73,70) := "11111111";
			tmp(73,71) := "11111111";
			tmp(73,72) := "11111111";
			tmp(73,73) := "11111111";
			tmp(73,74) := "11111111";
			tmp(73,75) := "11111111";
			tmp(73,76) := "11111111";
			tmp(73,77) := "11111111";
			tmp(73,78) := "11111111";
			tmp(73,79) := "11111111";
			tmp(73,80) := "11111111";
			tmp(74,1) := "11111111";
			tmp(74,2) := "11111111";
			tmp(74,3) := "11111111";
			tmp(74,4) := "11111111";
			tmp(74,5) := "11111111";
			tmp(74,6) := "11111111";
			tmp(74,7) := "11111111";
			tmp(74,8) := "11111111";
			tmp(74,9) := "11111111";
			tmp(74,10) := "11111111";
			tmp(74,11) := "11111111";
			tmp(74,12) := "11111111";
			tmp(74,13) := "11111111";
			tmp(74,14) := "11111111";
			tmp(74,15) := "11111111";
			tmp(74,16) := "11111111";
			tmp(74,17) := "11111111";
			tmp(74,18) := "11111111";
			tmp(74,19) := "11111101";
			tmp(74,20) := "11111111";
			tmp(74,21) := "11111111";
			tmp(74,22) := "11111111";
			tmp(74,23) := "11111111";
			tmp(74,24) := "11111100";
			tmp(74,25) := "11011111";
			tmp(74,26) := "11110011";
			tmp(74,27) := "11111111";
			tmp(74,28) := "11111111";
			tmp(74,29) := "11111111";
			tmp(74,30) := "11111100";
			tmp(74,31) := "11111010";
			tmp(74,32) := "11111101";
			tmp(74,33) := "11110111";
			tmp(74,34) := "11111111";
			tmp(74,35) := "11011010";
			tmp(74,36) := "01111011";
			tmp(74,37) := "11110111";
			tmp(74,38) := "11111101";
			tmp(74,39) := "11111111";
			tmp(74,40) := "11111100";
			tmp(74,41) := "11111000";
			tmp(74,42) := "11111011";
			tmp(74,43) := "11111101";
			tmp(74,44) := "11111111";
			tmp(74,45) := "11111111";
			tmp(74,46) := "11111110";
			tmp(74,47) := "11111111";
			tmp(74,48) := "11111111";
			tmp(74,49) := "11111111";
			tmp(74,50) := "11111111";
			tmp(74,51) := "11111111";
			tmp(74,52) := "11111111";
			tmp(74,53) := "11111111";
			tmp(74,54) := "11111111";
			tmp(74,55) := "11111111";
			tmp(74,56) := "11111111";
			tmp(74,57) := "11111111";
			tmp(74,58) := "11111111";
			tmp(74,59) := "11111111";
			tmp(74,60) := "11111111";
			tmp(74,61) := "11111111";
			tmp(74,62) := "11111111";
			tmp(74,63) := "11111111";
			tmp(74,64) := "11111111";
			tmp(74,65) := "11111111";
			tmp(74,66) := "11111111";
			tmp(74,67) := "11111111";
			tmp(74,68) := "11111111";
			tmp(74,69) := "11111111";
			tmp(74,70) := "11111111";
			tmp(74,71) := "11111111";
			tmp(74,72) := "11111111";
			tmp(74,73) := "11111111";
			tmp(74,74) := "11111111";
			tmp(74,75) := "11111111";
			tmp(74,76) := "11111111";
			tmp(74,77) := "11111111";
			tmp(74,78) := "11111111";
			tmp(74,79) := "11111111";
			tmp(74,80) := "11111111";
			tmp(75,1) := "11111111";
			tmp(75,2) := "11111111";
			tmp(75,3) := "11111111";
			tmp(75,4) := "11111111";
			tmp(75,5) := "11111111";
			tmp(75,6) := "11111111";
			tmp(75,7) := "11111111";
			tmp(75,8) := "11111111";
			tmp(75,9) := "11111111";
			tmp(75,10) := "11111111";
			tmp(75,11) := "11111111";
			tmp(75,12) := "11111111";
			tmp(75,13) := "11111111";
			tmp(75,14) := "11111111";
			tmp(75,15) := "11111111";
			tmp(75,16) := "11111111";
			tmp(75,17) := "11111110";
			tmp(75,18) := "11111111";
			tmp(75,19) := "11111111";
			tmp(75,20) := "11111111";
			tmp(75,21) := "11111111";
			tmp(75,22) := "11111111";
			tmp(75,23) := "11111111";
			tmp(75,24) := "11111111";
			tmp(75,25) := "11111101";
			tmp(75,26) := "11111111";
			tmp(75,27) := "11111111";
			tmp(75,28) := "11111110";
			tmp(75,29) := "11111111";
			tmp(75,30) := "11111111";
			tmp(75,31) := "11111110";
			tmp(75,32) := "11111111";
			tmp(75,33) := "11111100";
			tmp(75,34) := "11111110";
			tmp(75,35) := "10110001";
			tmp(75,36) := "10110110";
			tmp(75,37) := "11110101";
			tmp(75,38) := "11111111";
			tmp(75,39) := "11111110";
			tmp(75,40) := "11111111";
			tmp(75,41) := "11111110";
			tmp(75,42) := "11111101";
			tmp(75,43) := "11111110";
			tmp(75,44) := "11111111";
			tmp(75,45) := "11111110";
			tmp(75,46) := "11111110";
			tmp(75,47) := "11111111";
			tmp(75,48) := "11111110";
			tmp(75,49) := "11111111";
			tmp(75,50) := "11111111";
			tmp(75,51) := "11111111";
			tmp(75,52) := "11111111";
			tmp(75,53) := "11111111";
			tmp(75,54) := "11111111";
			tmp(75,55) := "11111111";
			tmp(75,56) := "11111111";
			tmp(75,57) := "11111111";
			tmp(75,58) := "11111111";
			tmp(75,59) := "11111111";
			tmp(75,60) := "11111111";
			tmp(75,61) := "11111111";
			tmp(75,62) := "11111111";
			tmp(75,63) := "11111111";
			tmp(75,64) := "11111111";
			tmp(75,65) := "11111111";
			tmp(75,66) := "11111111";
			tmp(75,67) := "11111111";
			tmp(75,68) := "11111111";
			tmp(75,69) := "11111111";
			tmp(75,70) := "11111111";
			tmp(75,71) := "11111111";
			tmp(75,72) := "11111111";
			tmp(75,73) := "11111111";
			tmp(75,74) := "11111111";
			tmp(75,75) := "11111111";
			tmp(75,76) := "11111111";
			tmp(75,77) := "11111111";
			tmp(75,78) := "11111111";
			tmp(75,79) := "11111111";
			tmp(75,80) := "11111111";
			tmp(76,1) := "11111111";
			tmp(76,2) := "11111111";
			tmp(76,3) := "11111111";
			tmp(76,4) := "11111111";
			tmp(76,5) := "11111111";
			tmp(76,6) := "11111111";
			tmp(76,7) := "11111111";
			tmp(76,8) := "11111111";
			tmp(76,9) := "11111111";
			tmp(76,10) := "11111111";
			tmp(76,11) := "11111111";
			tmp(76,12) := "11111111";
			tmp(76,13) := "11111111";
			tmp(76,14) := "11111111";
			tmp(76,15) := "11111111";
			tmp(76,16) := "11111111";
			tmp(76,17) := "11111111";
			tmp(76,18) := "11111111";
			tmp(76,19) := "11111111";
			tmp(76,20) := "11111110";
			tmp(76,21) := "11111110";
			tmp(76,22) := "11111111";
			tmp(76,23) := "11111111";
			tmp(76,24) := "11111101";
			tmp(76,25) := "11111100";
			tmp(76,26) := "11111100";
			tmp(76,27) := "11111110";
			tmp(76,28) := "11111100";
			tmp(76,29) := "11111010";
			tmp(76,30) := "11111110";
			tmp(76,31) := "11111110";
			tmp(76,32) := "11111100";
			tmp(76,33) := "11111110";
			tmp(76,34) := "11111101";
			tmp(76,35) := "11100101";
			tmp(76,36) := "11100000";
			tmp(76,37) := "11111110";
			tmp(76,38) := "11111111";
			tmp(76,39) := "11111111";
			tmp(76,40) := "11111111";
			tmp(76,41) := "11111101";
			tmp(76,42) := "11111111";
			tmp(76,43) := "11111111";
			tmp(76,44) := "11111110";
			tmp(76,45) := "11111110";
			tmp(76,46) := "11111111";
			tmp(76,47) := "11111111";
			tmp(76,48) := "11111110";
			tmp(76,49) := "11111111";
			tmp(76,50) := "11111111";
			tmp(76,51) := "11111111";
			tmp(76,52) := "11111111";
			tmp(76,53) := "11111111";
			tmp(76,54) := "11111111";
			tmp(76,55) := "11111111";
			tmp(76,56) := "11111111";
			tmp(76,57) := "11111111";
			tmp(76,58) := "11111111";
			tmp(76,59) := "11111111";
			tmp(76,60) := "11111111";
			tmp(76,61) := "11111111";
			tmp(76,62) := "11111111";
			tmp(76,63) := "11111111";
			tmp(76,64) := "11111111";
			tmp(76,65) := "11111111";
			tmp(76,66) := "11111111";
			tmp(76,67) := "11111111";
			tmp(76,68) := "11111111";
			tmp(76,69) := "11111111";
			tmp(76,70) := "11111111";
			tmp(76,71) := "11111111";
			tmp(76,72) := "11111111";
			tmp(76,73) := "11111111";
			tmp(76,74) := "11111111";
			tmp(76,75) := "11111111";
			tmp(76,76) := "11111111";
			tmp(76,77) := "11111111";
			tmp(76,78) := "11111111";
			tmp(76,79) := "11111111";
			tmp(76,80) := "11111111";
			tmp(77,1) := "11111111";
			tmp(77,2) := "11111111";
			tmp(77,3) := "11111111";
			tmp(77,4) := "11111111";
			tmp(77,5) := "11111111";
			tmp(77,6) := "11111111";
			tmp(77,7) := "11111111";
			tmp(77,8) := "11111111";
			tmp(77,9) := "11111111";
			tmp(77,10) := "11111111";
			tmp(77,11) := "11111111";
			tmp(77,12) := "11111111";
			tmp(77,13) := "11111111";
			tmp(77,14) := "11111111";
			tmp(77,15) := "11111111";
			tmp(77,16) := "11111111";
			tmp(77,17) := "11111111";
			tmp(77,18) := "11111101";
			tmp(77,19) := "11111111";
			tmp(77,20) := "11111111";
			tmp(77,21) := "11111110";
			tmp(77,22) := "11111111";
			tmp(77,23) := "11111111";
			tmp(77,24) := "11111111";
			tmp(77,25) := "11111110";
			tmp(77,26) := "11111111";
			tmp(77,27) := "11111110";
			tmp(77,28) := "11111111";
			tmp(77,29) := "11111110";
			tmp(77,30) := "11111111";
			tmp(77,31) := "11111111";
			tmp(77,32) := "11111111";
			tmp(77,33) := "11111111";
			tmp(77,34) := "11111111";
			tmp(77,35) := "11101100";
			tmp(77,36) := "11110110";
			tmp(77,37) := "11111110";
			tmp(77,38) := "11111111";
			tmp(77,39) := "11111110";
			tmp(77,40) := "11111111";
			tmp(77,41) := "11111111";
			tmp(77,42) := "11111111";
			tmp(77,43) := "11111111";
			tmp(77,44) := "11111110";
			tmp(77,45) := "11111111";
			tmp(77,46) := "11111111";
			tmp(77,47) := "11111110";
			tmp(77,48) := "11111111";
			tmp(77,49) := "11111111";
			tmp(77,50) := "11111111";
			tmp(77,51) := "11111111";
			tmp(77,52) := "11111111";
			tmp(77,53) := "11111111";
			tmp(77,54) := "11111111";
			tmp(77,55) := "11111111";
			tmp(77,56) := "11111111";
			tmp(77,57) := "11111111";
			tmp(77,58) := "11111111";
			tmp(77,59) := "11111111";
			tmp(77,60) := "11111111";
			tmp(77,61) := "11111111";
			tmp(77,62) := "11111111";
			tmp(77,63) := "11111111";
			tmp(77,64) := "11111111";
			tmp(77,65) := "11111111";
			tmp(77,66) := "11111111";
			tmp(77,67) := "11111111";
			tmp(77,68) := "11111111";
			tmp(77,69) := "11111111";
			tmp(77,70) := "11111111";
			tmp(77,71) := "11111111";
			tmp(77,72) := "11111111";
			tmp(77,73) := "11111111";
			tmp(77,74) := "11111111";
			tmp(77,75) := "11111111";
			tmp(77,76) := "11111111";
			tmp(77,77) := "11111111";
			tmp(77,78) := "11111111";
			tmp(77,79) := "11111111";
			tmp(77,80) := "11111111";
			tmp(78,1) := "11111111";
			tmp(78,2) := "11111111";
			tmp(78,3) := "11111111";
			tmp(78,4) := "11111111";
			tmp(78,5) := "11111111";
			tmp(78,6) := "11111111";
			tmp(78,7) := "11111111";
			tmp(78,8) := "11111111";
			tmp(78,9) := "11111111";
			tmp(78,10) := "11111111";
			tmp(78,11) := "11111111";
			tmp(78,12) := "11111111";
			tmp(78,13) := "11111111";
			tmp(78,14) := "11111111";
			tmp(78,15) := "11111111";
			tmp(78,16) := "11111111";
			tmp(78,17) := "11111111";
			tmp(78,18) := "11111110";
			tmp(78,19) := "11111111";
			tmp(78,20) := "11111111";
			tmp(78,21) := "11111111";
			tmp(78,22) := "11111111";
			tmp(78,23) := "11111101";
			tmp(78,24) := "11111111";
			tmp(78,25) := "11111111";
			tmp(78,26) := "11111110";
			tmp(78,27) := "11111111";
			tmp(78,28) := "11111111";
			tmp(78,29) := "11111111";
			tmp(78,30) := "11111111";
			tmp(78,31) := "11111110";
			tmp(78,32) := "11111111";
			tmp(78,33) := "11111111";
			tmp(78,34) := "11111111";
			tmp(78,35) := "11111101";
			tmp(78,36) := "11111111";
			tmp(78,37) := "11111011";
			tmp(78,38) := "11111111";
			tmp(78,39) := "11111110";
			tmp(78,40) := "11111110";
			tmp(78,41) := "11111111";
			tmp(78,42) := "11111110";
			tmp(78,43) := "11111111";
			tmp(78,44) := "11111111";
			tmp(78,45) := "11111111";
			tmp(78,46) := "11111111";
			tmp(78,47) := "11111110";
			tmp(78,48) := "11111111";
			tmp(78,49) := "11111111";
			tmp(78,50) := "11111111";
			tmp(78,51) := "11111111";
			tmp(78,52) := "11111111";
			tmp(78,53) := "11111111";
			tmp(78,54) := "11111111";
			tmp(78,55) := "11111111";
			tmp(78,56) := "11111111";
			tmp(78,57) := "11111111";
			tmp(78,58) := "11111111";
			tmp(78,59) := "11111111";
			tmp(78,60) := "11111111";
			tmp(78,61) := "11111111";
			tmp(78,62) := "11111111";
			tmp(78,63) := "11111111";
			tmp(78,64) := "11111111";
			tmp(78,65) := "11111111";
			tmp(78,66) := "11111111";
			tmp(78,67) := "11111111";
			tmp(78,68) := "11111111";
			tmp(78,69) := "11111111";
			tmp(78,70) := "11111111";
			tmp(78,71) := "11111111";
			tmp(78,72) := "11111111";
			tmp(78,73) := "11111111";
			tmp(78,74) := "11111111";
			tmp(78,75) := "11111111";
			tmp(78,76) := "11111111";
			tmp(78,77) := "11111111";
			tmp(78,78) := "11111111";
			tmp(78,79) := "11111111";
			tmp(78,80) := "11111111";
			tmp(79,1) := "11111111";
			tmp(79,2) := "11111111";
			tmp(79,3) := "11111111";
			tmp(79,4) := "11111111";
			tmp(79,5) := "11111111";
			tmp(79,6) := "11111111";
			tmp(79,7) := "11111111";
			tmp(79,8) := "11111111";
			tmp(79,9) := "11111111";
			tmp(79,10) := "11111111";
			tmp(79,11) := "11111111";
			tmp(79,12) := "11111111";
			tmp(79,13) := "11111111";
			tmp(79,14) := "11111111";
			tmp(79,15) := "11111111";
			tmp(79,16) := "11111111";
			tmp(79,17) := "11111111";
			tmp(79,18) := "11111111";
			tmp(79,19) := "11111110";
			tmp(79,20) := "11111110";
			tmp(79,21) := "11111111";
			tmp(79,22) := "11111111";
			tmp(79,23) := "11111111";
			tmp(79,24) := "11111111";
			tmp(79,25) := "11111111";
			tmp(79,26) := "11111110";
			tmp(79,27) := "11111100";
			tmp(79,28) := "11111110";
			tmp(79,29) := "11111110";
			tmp(79,30) := "11111110";
			tmp(79,31) := "11111110";
			tmp(79,32) := "11111100";
			tmp(79,33) := "11111110";
			tmp(79,34) := "11111111";
			tmp(79,35) := "11111101";
			tmp(79,36) := "11111111";
			tmp(79,37) := "11111110";
			tmp(79,38) := "11111111";
			tmp(79,39) := "11111101";
			tmp(79,40) := "11111111";
			tmp(79,41) := "11111110";
			tmp(79,42) := "11111111";
			tmp(79,43) := "11111111";
			tmp(79,44) := "11111111";
			tmp(79,45) := "11111110";
			tmp(79,46) := "11111111";
			tmp(79,47) := "11111111";
			tmp(79,48) := "11111111";
			tmp(79,49) := "11111111";
			tmp(79,50) := "11111111";
			tmp(79,51) := "11111111";
			tmp(79,52) := "11111111";
			tmp(79,53) := "11111111";
			tmp(79,54) := "11111111";
			tmp(79,55) := "11111111";
			tmp(79,56) := "11111111";
			tmp(79,57) := "11111111";
			tmp(79,58) := "11111111";
			tmp(79,59) := "11111111";
			tmp(79,60) := "11111111";
			tmp(79,61) := "11111111";
			tmp(79,62) := "11111111";
			tmp(79,63) := "11111111";
			tmp(79,64) := "11111111";
			tmp(79,65) := "11111111";
			tmp(79,66) := "11111111";
			tmp(79,67) := "11111111";
			tmp(79,68) := "11111111";
			tmp(79,69) := "11111111";
			tmp(79,70) := "11111111";
			tmp(79,71) := "11111111";
			tmp(79,72) := "11111111";
			tmp(79,73) := "11111111";
			tmp(79,74) := "11111111";
			tmp(79,75) := "11111111";
			tmp(79,76) := "11111111";
			tmp(79,77) := "11111111";
			tmp(79,78) := "11111111";
			tmp(79,79) := "11111111";
			tmp(79,80) := "11111111";
			tmp(80,1) := "11111111";
			tmp(80,2) := "11111111";
			tmp(80,3) := "11111111";
			tmp(80,4) := "11111111";
			tmp(80,5) := "11111111";
			tmp(80,6) := "11111111";
			tmp(80,7) := "11111111";
			tmp(80,8) := "11111111";
			tmp(80,9) := "11111111";
			tmp(80,10) := "11111111";
			tmp(80,11) := "11111111";
			tmp(80,12) := "11111111";
			tmp(80,13) := "11111111";
			tmp(80,14) := "11111111";
			tmp(80,15) := "11111111";
			tmp(80,16) := "11111111";
			tmp(80,17) := "11111111";
			tmp(80,18) := "11111111";
			tmp(80,19) := "11111110";
			tmp(80,20) := "11111111";
			tmp(80,21) := "11111111";
			tmp(80,22) := "11111110";
			tmp(80,23) := "11111111";
			tmp(80,24) := "11111111";
			tmp(80,25) := "11111111";
			tmp(80,26) := "11111111";
			tmp(80,27) := "11111110";
			tmp(80,28) := "11111110";
			tmp(80,29) := "11111111";
			tmp(80,30) := "11111111";
			tmp(80,31) := "11111111";
			tmp(80,32) := "11111100";
			tmp(80,33) := "11111110";
			tmp(80,34) := "11111101";
			tmp(80,35) := "11111100";
			tmp(80,36) := "11111111";
			tmp(80,37) := "11111110";
			tmp(80,38) := "11111110";
			tmp(80,39) := "11111110";
			tmp(80,40) := "11111111";
			tmp(80,41) := "11111111";
			tmp(80,42) := "11111111";
			tmp(80,43) := "11111110";
			tmp(80,44) := "11111101";
			tmp(80,45) := "11111111";
			tmp(80,46) := "11111111";
			tmp(80,47) := "11111110";
			tmp(80,48) := "11111111";
			tmp(80,49) := "11111111";
			tmp(80,50) := "11111111";
			tmp(80,51) := "11111111";
			tmp(80,52) := "11111111";
			tmp(80,53) := "11111111";
			tmp(80,54) := "11111111";
			tmp(80,55) := "11111111";
			tmp(80,56) := "11111111";
			tmp(80,57) := "11111111";
			tmp(80,58) := "11111111";
			tmp(80,59) := "11111111";
			tmp(80,60) := "11111111";
			tmp(80,61) := "11111111";
			tmp(80,62) := "11111111";
			tmp(80,63) := "11111111";
			tmp(80,64) := "11111111";
			tmp(80,65) := "11111111";
			tmp(80,66) := "11111111";
			tmp(80,67) := "11111111";
			tmp(80,68) := "11111111";
			tmp(80,69) := "11111111";
			tmp(80,70) := "11111111";
			tmp(80,71) := "11111111";
			tmp(80,72) := "11111111";
			tmp(80,73) := "11111111";
			tmp(80,74) := "11111111";
			tmp(80,75) := "11111111";
			tmp(80,76) := "11111111";
			tmp(80,77) := "11111111";
			tmp(80,78) := "11111111";
			tmp(80,79) := "11111111";
			tmp(80,80) := "11111111";

		return tmp;
	end init_rom;
	
	-- Declare the ROM signal and specify a default value.	Quartus II
	-- will create a memory initialization file (.mif) based on the 
	-- default value.
	signal rom : memory_t := init_rom;
begin
	process(clk)
	variable t : matrix_in;
	begin
		for i in addr_i to (addr_i + elin-1) loop
			for j in addr_j to (addr_j + ecol-1) loop
				t(i, j) := rom(addr_i+i, addr_j+j);
			end loop;
		end loop;
		if(rising_edge(clk)) then
			q <= t;
		end if;
	end process;
		
end rtl;
