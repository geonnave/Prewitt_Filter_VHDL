library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package mem_size is
	constant	col	:	integer	:=	38;			-->	
	constant	lin	:	integer	:=	38;			-->	
end;
